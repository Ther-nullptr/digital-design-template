//$Id: xor.genpp,v 1.5 2006/06/13 06:30:06 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module XOR3X4MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  xor I0(Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
     if ((B == 1'b1) && (C == 1'b1))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b1) && (C == 1'b0))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b0) && (C == 1'b1))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b0) && (C == 1'b0))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((A == 1'b1) && (C == 1'b1))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b1) && (C == 1'b0))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b0) && (C == 1'b1))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b0) && (C == 1'b0))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
    if (A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify

endmodule // XOR3X4MA10TR
`endcelldefine
//$Id: xor.genpp,v 1.5 2006/06/13 06:30:06 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module XOR3X3MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  xor I0(Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
     if ((B == 1'b1) && (C == 1'b1))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b1) && (C == 1'b0))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b0) && (C == 1'b1))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b0) && (C == 1'b0))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((A == 1'b1) && (C == 1'b1))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b1) && (C == 1'b0))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b0) && (C == 1'b1))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b0) && (C == 1'b0))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
    if (A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify

endmodule // XOR3X3MA10TR
`endcelldefine
//$Id: xor.genpp,v 1.5 2006/06/13 06:30:06 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module XOR3X2MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  xor I0(Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
     if ((B == 1'b1) && (C == 1'b1))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b1) && (C == 1'b0))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b0) && (C == 1'b1))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b0) && (C == 1'b0))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((A == 1'b1) && (C == 1'b1))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b1) && (C == 1'b0))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b0) && (C == 1'b1))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b0) && (C == 1'b0))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
    if (A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify

endmodule // XOR3X2MA10TR
`endcelldefine
//$Id: xor.genpp,v 1.5 2006/06/13 06:30:06 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module XOR3X1P4MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  xor I0(Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
     if ((B == 1'b1) && (C == 1'b1))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b1) && (C == 1'b0))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b0) && (C == 1'b1))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b0) && (C == 1'b0))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((A == 1'b1) && (C == 1'b1))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b1) && (C == 1'b0))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b0) && (C == 1'b1))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b0) && (C == 1'b0))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
    if (A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify

endmodule // XOR3X1P4MA10TR
`endcelldefine
//$Id: xor.genpp,v 1.5 2006/06/13 06:30:06 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module XOR3X1MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  xor I0(Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
     if ((B == 1'b1) && (C == 1'b1))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b1) && (C == 1'b0))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b0) && (C == 1'b1))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b0) && (C == 1'b0))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((A == 1'b1) && (C == 1'b1))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b1) && (C == 1'b0))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b0) && (C == 1'b1))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b0) && (C == 1'b0))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
    if (A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify

endmodule // XOR3X1MA10TR
`endcelldefine
//$Id: xor.genpp,v 1.5 2006/06/13 06:30:06 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module XOR3X0P7MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  xor I0(Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
     if ((B == 1'b1) && (C == 1'b1))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b1) && (C == 1'b0))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b0) && (C == 1'b1))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b0) && (C == 1'b0))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((A == 1'b1) && (C == 1'b1))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b1) && (C == 1'b0))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b0) && (C == 1'b1))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b0) && (C == 1'b0))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
    if (A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify

endmodule // XOR3X0P7MA10TR
`endcelldefine
//$Id: xor.genpp,v 1.5 2006/06/13 06:30:06 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module XOR3X0P5MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  xor I0(Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
     if ((B == 1'b1) && (C == 1'b1))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b1) && (C == 1'b0))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b0) && (C == 1'b1))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b0) && (C == 1'b0))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((A == 1'b1) && (C == 1'b1))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b1) && (C == 1'b0))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b0) && (C == 1'b1))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b0) && (C == 1'b0))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
    if (A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify

endmodule // XOR3X0P5MA10TR
`endcelldefine
//$Id: xor.genpp,v 1.5 2006/06/13 06:30:06 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module XOR2X4MA10TR (Y, A, B);
output Y;
input A, B;

  xor I0(Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
     if (B == 1'b1)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (B == 1'b0)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (A == 1'b1)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if (A == 1'b0)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // XOR2X4MA10TR
`endcelldefine
//$Id: xor.genpp,v 1.5 2006/06/13 06:30:06 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module XOR2X3MA10TR (Y, A, B);
output Y;
input A, B;

  xor I0(Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
     if (B == 1'b1)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (B == 1'b0)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (A == 1'b1)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if (A == 1'b0)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // XOR2X3MA10TR
`endcelldefine
//$Id: xor.genpp,v 1.5 2006/06/13 06:30:06 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module XOR2X2MA10TR (Y, A, B);
output Y;
input A, B;

  xor I0(Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
     if (B == 1'b1)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (B == 1'b0)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (A == 1'b1)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if (A == 1'b0)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // XOR2X2MA10TR
`endcelldefine
//$Id: xor.genpp,v 1.5 2006/06/13 06:30:06 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module XOR2X1P4MA10TR (Y, A, B);
output Y;
input A, B;

  xor I0(Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
     if (B == 1'b1)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (B == 1'b0)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (A == 1'b1)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if (A == 1'b0)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // XOR2X1P4MA10TR
`endcelldefine
//$Id: xor.genpp,v 1.5 2006/06/13 06:30:06 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module XOR2X1MA10TR (Y, A, B);
output Y;
input A, B;

  xor I0(Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
     if (B == 1'b1)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (B == 1'b0)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (A == 1'b1)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if (A == 1'b0)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // XOR2X1MA10TR
`endcelldefine
//$Id: xor.genpp,v 1.5 2006/06/13 06:30:06 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module XOR2X0P7MA10TR (Y, A, B);
output Y;
input A, B;

  xor I0(Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
     if (B == 1'b1)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (B == 1'b0)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (A == 1'b1)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if (A == 1'b0)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // XOR2X0P7MA10TR
`endcelldefine
//$Id: xor.genpp,v 1.5 2006/06/13 06:30:06 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module XOR2X0P5MA10TR (Y, A, B);
output Y;
input A, B;

  xor I0(Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
     if (B == 1'b1)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (B == 1'b0)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (A == 1'b1)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if (A == 1'b0)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // XOR2X0P5MA10TR
`endcelldefine
//$Id: xor.genpp,v 1.5 2006/06/13 06:30:06 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module XNOR3X4MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  xnor I0(Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
     if ((B == 1'b1) && (C == 1'b1))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b1) && (C == 1'b0))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b0) && (C == 1'b1))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b0) && (C == 1'b0))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((A == 1'b1) && (C == 1'b1))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b1) && (C == 1'b0))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b0) && (C == 1'b1))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b0) && (C == 1'b0))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
    if (A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify

endmodule // XNOR3X4MA10TR
`endcelldefine
//$Id: xor.genpp,v 1.5 2006/06/13 06:30:06 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module XNOR3X3MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  xnor I0(Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
     if ((B == 1'b1) && (C == 1'b1))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b1) && (C == 1'b0))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b0) && (C == 1'b1))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b0) && (C == 1'b0))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((A == 1'b1) && (C == 1'b1))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b1) && (C == 1'b0))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b0) && (C == 1'b1))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b0) && (C == 1'b0))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
    if (A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify

endmodule // XNOR3X3MA10TR
`endcelldefine
//$Id: xor.genpp,v 1.5 2006/06/13 06:30:06 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module XNOR3X2MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  xnor I0(Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
     if ((B == 1'b1) && (C == 1'b1))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b1) && (C == 1'b0))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b0) && (C == 1'b1))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b0) && (C == 1'b0))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((A == 1'b1) && (C == 1'b1))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b1) && (C == 1'b0))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b0) && (C == 1'b1))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b0) && (C == 1'b0))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
    if (A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify

endmodule // XNOR3X2MA10TR
`endcelldefine
//$Id: xor.genpp,v 1.5 2006/06/13 06:30:06 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module XNOR3X1P4MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  xnor I0(Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
     if ((B == 1'b1) && (C == 1'b1))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b1) && (C == 1'b0))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b0) && (C == 1'b1))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b0) && (C == 1'b0))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((A == 1'b1) && (C == 1'b1))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b1) && (C == 1'b0))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b0) && (C == 1'b1))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b0) && (C == 1'b0))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
    if (A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify

endmodule // XNOR3X1P4MA10TR
`endcelldefine
//$Id: xor.genpp,v 1.5 2006/06/13 06:30:06 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module XNOR3X1MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  xnor I0(Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
     if ((B == 1'b1) && (C == 1'b1))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b1) && (C == 1'b0))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b0) && (C == 1'b1))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b0) && (C == 1'b0))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((A == 1'b1) && (C == 1'b1))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b1) && (C == 1'b0))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b0) && (C == 1'b1))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b0) && (C == 1'b0))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
    if (A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify

endmodule // XNOR3X1MA10TR
`endcelldefine
//$Id: xor.genpp,v 1.5 2006/06/13 06:30:06 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module XNOR3X0P7MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  xnor I0(Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
     if ((B == 1'b1) && (C == 1'b1))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b1) && (C == 1'b0))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b0) && (C == 1'b1))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b0) && (C == 1'b0))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((A == 1'b1) && (C == 1'b1))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b1) && (C == 1'b0))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b0) && (C == 1'b1))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b0) && (C == 1'b0))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
    if (A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify

endmodule // XNOR3X0P7MA10TR
`endcelldefine
//$Id: xor.genpp,v 1.5 2006/06/13 06:30:06 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module XNOR3X0P5MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  xnor I0(Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
     if ((B == 1'b1) && (C == 1'b1))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b1) && (C == 1'b0))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b0) && (C == 1'b1))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((B == 1'b0) && (C == 1'b0))
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if ((A == 1'b1) && (C == 1'b1))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b1) && (C == 1'b0))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b0) && (C == 1'b1))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if ((A == 1'b0) && (C == 1'b0))
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
    if (A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify

endmodule // XNOR3X0P5MA10TR
`endcelldefine
//$Id: xor.genpp,v 1.5 2006/06/13 06:30:06 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module XNOR2X4MA10TR (Y, A, B);
output Y;
input A, B;

  xnor I0(Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
     if (B == 1'b1)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (B == 1'b0)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (A == 1'b1)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if (A == 1'b0)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // XNOR2X4MA10TR
`endcelldefine
//$Id: xor.genpp,v 1.5 2006/06/13 06:30:06 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module XNOR2X3MA10TR (Y, A, B);
output Y;
input A, B;

  xnor I0(Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
     if (B == 1'b1)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (B == 1'b0)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (A == 1'b1)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if (A == 1'b0)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // XNOR2X3MA10TR
`endcelldefine
//$Id: xor.genpp,v 1.5 2006/06/13 06:30:06 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module XNOR2X2MA10TR (Y, A, B);
output Y;
input A, B;

  xnor I0(Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
     if (B == 1'b1)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (B == 1'b0)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (A == 1'b1)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if (A == 1'b0)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // XNOR2X2MA10TR
`endcelldefine
//$Id: xor.genpp,v 1.5 2006/06/13 06:30:06 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module XNOR2X1P4MA10TR (Y, A, B);
output Y;
input A, B;

  xnor I0(Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
     if (B == 1'b1)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (B == 1'b0)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (A == 1'b1)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if (A == 1'b0)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // XNOR2X1P4MA10TR
`endcelldefine
//$Id: xor.genpp,v 1.5 2006/06/13 06:30:06 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module XNOR2X1MA10TR (Y, A, B);
output Y;
input A, B;

  xnor I0(Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
     if (B == 1'b1)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (B == 1'b0)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (A == 1'b1)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if (A == 1'b0)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // XNOR2X1MA10TR
`endcelldefine
//$Id: xor.genpp,v 1.5 2006/06/13 06:30:06 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module XNOR2X0P7MA10TR (Y, A, B);
output Y;
input A, B;

  xnor I0(Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
     if (B == 1'b1)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (B == 1'b0)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (A == 1'b1)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if (A == 1'b0)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // XNOR2X0P7MA10TR
`endcelldefine
//$Id: xor.genpp,v 1.5 2006/06/13 06:30:06 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module XNOR2X0P5MA10TR (Y, A, B);
output Y;
input A, B;

  xnor I0(Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
     if (B == 1'b1)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (B == 1'b0)
	(A *> Y) = (tplh$A$Y, tphl$A$Y);
     if (A == 1'b1)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
     if (A == 1'b0)
	(B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // XNOR2X0P5MA10TR
`endcelldefine
//$Id: tie.genpp,v 1.1.1.1 2002/12/05 17:56:00 ron Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module TIELOX1MA10TR (Y);
output Y;

  buf I0(Y, 1'b0);

endmodule //TIELOX1MA10TR 
`endcelldefine
//$Id: tie.genpp,v 1.1.1.1 2002/12/05 17:56:00 ron Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module TIEHIX1MA10TR (Y);
output Y;

  buf I0(Y, 1'b1);

endmodule //TIEHIX1MA10TR 
`endcelldefine
//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFYQX4MA10TR (Q, D, SI, SE, CK);
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // SDFFYQX4MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFYQX3MA10TR (Q, D, SI, SE, CK);
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // SDFFYQX3MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFYQX2MA10TR (Q, D, SI, SE, CK);
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // SDFFYQX2MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFYQX1MA10TR (Q, D, SI, SE, CK);
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // SDFFYQX1MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFSRPQX4MA10TR (Q, D, SI, SE, CK, SN, R);
output Q;
input D, SI, SE, CK, SN, R;
reg NOTIFIER;
  not   XX0 (xRN, R);
  buf   XX1 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$SN$Q = 1.0,
      tphl$SN$Q = 1.0,
      tplh$R$Q = 1.0,
      tphl$R$Q = 1.0,
      tminpwl$SN = 1.0,
      tminpwh$SN = 1.0,
      tminpwl$R = 1.0,
      tminpwh$R = 1.0,
      tsetup$SN$CK = 1.0,
      thold$SN$CK = 0.5,
      tsetup$R$CK = 1.0,
      thold$R$CK = 0.5,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      thold$R$SN = 1.0,
      thold$SN$R = 1.0,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK, negedge R &&& (SN == 1'b1), tsetup$R$CK ,thold$R$CK , NOTIFIER);
    $width(posedge R &&& (SN == 1'b1), tminpwh$R, 0, NOTIFIER);
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK ,thold$SN$CK , NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    $hold(negedge R, negedge SN, thold$SN$R, NOTIFIER);    
    $hold(posedge SN, posedge R, thold$R$SN, NOTIFIER);    
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 

endspecify
endmodule // SDFFSRPQX4MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFSRPQX3MA10TR (Q, D, SI, SE, CK, SN, R);
output Q;
input D, SI, SE, CK, SN, R;
reg NOTIFIER;
  not   XX0 (xRN, R);
  buf   XX1 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$SN$Q = 1.0,
      tphl$SN$Q = 1.0,
      tplh$R$Q = 1.0,
      tphl$R$Q = 1.0,
      tminpwl$SN = 1.0,
      tminpwh$SN = 1.0,
      tminpwl$R = 1.0,
      tminpwh$R = 1.0,
      tsetup$SN$CK = 1.0,
      thold$SN$CK = 0.5,
      tsetup$R$CK = 1.0,
      thold$R$CK = 0.5,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      thold$R$SN = 1.0,
      thold$SN$R = 1.0,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK, negedge R &&& (SN == 1'b1), tsetup$R$CK ,thold$R$CK , NOTIFIER);
    $width(posedge R &&& (SN == 1'b1), tminpwh$R, 0, NOTIFIER);
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK ,thold$SN$CK , NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    $hold(negedge R, negedge SN, thold$SN$R, NOTIFIER);    
    $hold(posedge SN, posedge R, thold$R$SN, NOTIFIER);    
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 

endspecify
endmodule // SDFFSRPQX3MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFSRPQX2MA10TR (Q, D, SI, SE, CK, SN, R);
output Q;
input D, SI, SE, CK, SN, R;
reg NOTIFIER;
  not   XX0 (xRN, R);
  buf   XX1 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$SN$Q = 1.0,
      tphl$SN$Q = 1.0,
      tplh$R$Q = 1.0,
      tphl$R$Q = 1.0,
      tminpwl$SN = 1.0,
      tminpwh$SN = 1.0,
      tminpwl$R = 1.0,
      tminpwh$R = 1.0,
      tsetup$SN$CK = 1.0,
      thold$SN$CK = 0.5,
      tsetup$R$CK = 1.0,
      thold$R$CK = 0.5,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      thold$R$SN = 1.0,
      thold$SN$R = 1.0,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK, negedge R &&& (SN == 1'b1), tsetup$R$CK ,thold$R$CK , NOTIFIER);
    $width(posedge R &&& (SN == 1'b1), tminpwh$R, 0, NOTIFIER);
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK ,thold$SN$CK , NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    $hold(negedge R, negedge SN, thold$SN$R, NOTIFIER);    
    $hold(posedge SN, posedge R, thold$R$SN, NOTIFIER);    
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 

endspecify
endmodule // SDFFSRPQX2MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFSRPQX1MA10TR (Q, D, SI, SE, CK, SN, R);
output Q;
input D, SI, SE, CK, SN, R;
reg NOTIFIER;
  not   XX0 (xRN, R);
  buf   XX1 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$SN$Q = 1.0,
      tphl$SN$Q = 1.0,
      tplh$R$Q = 1.0,
      tphl$R$Q = 1.0,
      tminpwl$SN = 1.0,
      tminpwh$SN = 1.0,
      tminpwl$R = 1.0,
      tminpwh$R = 1.0,
      tsetup$SN$CK = 1.0,
      thold$SN$CK = 0.5,
      tsetup$R$CK = 1.0,
      thold$R$CK = 0.5,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      thold$R$SN = 1.0,
      thold$SN$R = 1.0,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK, negedge R &&& (SN == 1'b1), tsetup$R$CK ,thold$R$CK , NOTIFIER);
    $width(posedge R &&& (SN == 1'b1), tminpwh$R, 0, NOTIFIER);
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK ,thold$SN$CK , NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    $hold(negedge R, negedge SN, thold$SN$R, NOTIFIER);    
    $hold(posedge SN, posedge R, thold$R$SN, NOTIFIER);    
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 

endspecify
endmodule // SDFFSRPQX1MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFSRPQX0P5MA10TR (Q, D, SI, SE, CK, SN, R);
output Q;
input D, SI, SE, CK, SN, R;
reg NOTIFIER;
  not   XX0 (xRN, R);
  buf   XX1 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$SN$Q = 1.0,
      tphl$SN$Q = 1.0,
      tplh$R$Q = 1.0,
      tphl$R$Q = 1.0,
      tminpwl$SN = 1.0,
      tminpwh$SN = 1.0,
      tminpwl$R = 1.0,
      tminpwh$R = 1.0,
      tsetup$SN$CK = 1.0,
      thold$SN$CK = 0.5,
      tsetup$R$CK = 1.0,
      thold$R$CK = 0.5,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      thold$R$SN = 1.0,
      thold$SN$R = 1.0,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK, negedge R &&& (SN == 1'b1), tsetup$R$CK ,thold$R$CK , NOTIFIER);
    $width(posedge R &&& (SN == 1'b1), tminpwh$R, 0, NOTIFIER);
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK ,thold$SN$CK , NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    $hold(negedge R, negedge SN, thold$SN$R, NOTIFIER);    
    $hold(posedge SN, posedge R, thold$R$SN, NOTIFIER);    
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 

endspecify
endmodule // SDFFSRPQX0P5MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFSQNX3MA10TR (QN, D, SI, SE, CK, SN);
output QN;
input D, SI, SE, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  not     I72 (QN, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$SN$QN = 1.0,
      tphl$SN$QN = 1.0,
      tminpwl$SN = 1.0,
      tminpwh$SN = 1.0,
      tsetup$SN$CK = 1.0,
      thold$SN$CK = 0.5,
      tplh$CK$QN = 1.0,
      tphl$CK$QN = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (QN -: D)) = (tplh$CK$QN, tphl$CK$QN);
    if ( SandRandSE )
      (posedge CK *> (QN -: SI)) = (tplh$CK$QN, tphl$CK$QN);

// timing checks
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK ,thold$SN$CK , NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 

endspecify
endmodule // SDFFSQNX3MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFSQNX2MA10TR (QN, D, SI, SE, CK, SN);
output QN;
input D, SI, SE, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  not     I72 (QN, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$SN$QN = 1.0,
      tphl$SN$QN = 1.0,
      tminpwl$SN = 1.0,
      tminpwh$SN = 1.0,
      tsetup$SN$CK = 1.0,
      thold$SN$CK = 0.5,
      tplh$CK$QN = 1.0,
      tphl$CK$QN = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (QN -: D)) = (tplh$CK$QN, tphl$CK$QN);
    if ( SandRandSE )
      (posedge CK *> (QN -: SI)) = (tplh$CK$QN, tphl$CK$QN);

// timing checks
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK ,thold$SN$CK , NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 

endspecify
endmodule // SDFFSQNX2MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFSQNX1MA10TR (QN, D, SI, SE, CK, SN);
output QN;
input D, SI, SE, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  not     I72 (QN, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$SN$QN = 1.0,
      tphl$SN$QN = 1.0,
      tminpwl$SN = 1.0,
      tminpwh$SN = 1.0,
      tsetup$SN$CK = 1.0,
      thold$SN$CK = 0.5,
      tplh$CK$QN = 1.0,
      tphl$CK$QN = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (QN -: D)) = (tplh$CK$QN, tphl$CK$QN);
    if ( SandRandSE )
      (posedge CK *> (QN -: SI)) = (tplh$CK$QN, tphl$CK$QN);

// timing checks
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK ,thold$SN$CK , NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 

endspecify
endmodule // SDFFSQNX1MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFSQNX0P5MA10TR (QN, D, SI, SE, CK, SN);
output QN;
input D, SI, SE, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  not     I72 (QN, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$SN$QN = 1.0,
      tphl$SN$QN = 1.0,
      tminpwl$SN = 1.0,
      tminpwh$SN = 1.0,
      tsetup$SN$CK = 1.0,
      thold$SN$CK = 0.5,
      tplh$CK$QN = 1.0,
      tphl$CK$QN = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (QN -: D)) = (tplh$CK$QN, tphl$CK$QN);
    if ( SandRandSE )
      (posedge CK *> (QN -: SI)) = (tplh$CK$QN, tphl$CK$QN);

// timing checks
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK ,thold$SN$CK , NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tphl$SN$QN); 

endspecify
endmodule // SDFFSQNX0P5MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFSQX4MA10TR (Q, D, SI, SE, CK, SN);
output Q;
input D, SI, SE, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$SN$Q = 1.0,
      tphl$SN$Q = 1.0,
      tminpwl$SN = 1.0,
      tminpwh$SN = 1.0,
      tsetup$SN$CK = 1.0,
      thold$SN$CK = 0.5,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK ,thold$SN$CK , NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q);

endspecify
endmodule // SDFFSQX4MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFSQX3MA10TR (Q, D, SI, SE, CK, SN);
output Q;
input D, SI, SE, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$SN$Q = 1.0,
      tphl$SN$Q = 1.0,
      tminpwl$SN = 1.0,
      tminpwh$SN = 1.0,
      tsetup$SN$CK = 1.0,
      thold$SN$CK = 0.5,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK ,thold$SN$CK , NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q);

endspecify
endmodule // SDFFSQX3MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFSQX2MA10TR (Q, D, SI, SE, CK, SN);
output Q;
input D, SI, SE, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$SN$Q = 1.0,
      tphl$SN$Q = 1.0,
      tminpwl$SN = 1.0,
      tminpwh$SN = 1.0,
      tsetup$SN$CK = 1.0,
      thold$SN$CK = 0.5,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK ,thold$SN$CK , NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q);

endspecify
endmodule // SDFFSQX2MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFSQX1MA10TR (Q, D, SI, SE, CK, SN);
output Q;
input D, SI, SE, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$SN$Q = 1.0,
      tphl$SN$Q = 1.0,
      tminpwl$SN = 1.0,
      tminpwh$SN = 1.0,
      tsetup$SN$CK = 1.0,
      thold$SN$CK = 0.5,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK ,thold$SN$CK , NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q);

endspecify
endmodule // SDFFSQX1MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFSQX0P5MA10TR (Q, D, SI, SE, CK, SN);
output Q;
input D, SI, SE, CK, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$SN$Q = 1.0,
      tphl$SN$Q = 1.0,
      tminpwl$SN = 1.0,
      tminpwh$SN = 1.0,
      tsetup$SN$CK = 1.0,
      thold$SN$CK = 0.5,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK ,thold$SN$CK , NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q);

endspecify
endmodule // SDFFSQX0P5MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFRPQNX3MA10TR (QN, D, SI, SE, CK, R);
output QN;
input D, SI, SE, CK, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  not     I72 (QN, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$R$QN = 1.0,
      tphl$R$QN = 1.0,
      tminpwl$R = 1.0,
      tminpwh$R = 1.0,
      tsetup$R$CK = 1.0,
      thold$R$CK = 0.5,
      tplh$CK$QN = 1.0,
      tphl$CK$QN = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (QN -: D)) = (tplh$CK$QN, tphl$CK$QN);
    if ( SandRandSE )
      (posedge CK *> (QN -: SI)) = (tplh$CK$QN, tphl$CK$QN);

// timing checks
    $setuphold(posedge CK, negedge R, tsetup$R$CK ,thold$R$CK , NOTIFIER);
    $width(posedge R, tminpwh$R, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 

endspecify
endmodule // SDFFRPQNX3MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFRPQNX2MA10TR (QN, D, SI, SE, CK, R);
output QN;
input D, SI, SE, CK, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  not     I72 (QN, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$R$QN = 1.0,
      tphl$R$QN = 1.0,
      tminpwl$R = 1.0,
      tminpwh$R = 1.0,
      tsetup$R$CK = 1.0,
      thold$R$CK = 0.5,
      tplh$CK$QN = 1.0,
      tphl$CK$QN = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (QN -: D)) = (tplh$CK$QN, tphl$CK$QN);
    if ( SandRandSE )
      (posedge CK *> (QN -: SI)) = (tplh$CK$QN, tphl$CK$QN);

// timing checks
    $setuphold(posedge CK, negedge R, tsetup$R$CK ,thold$R$CK , NOTIFIER);
    $width(posedge R, tminpwh$R, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 

endspecify
endmodule // SDFFRPQNX2MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFRPQNX1MA10TR (QN, D, SI, SE, CK, R);
output QN;
input D, SI, SE, CK, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  not     I72 (QN, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$R$QN = 1.0,
      tphl$R$QN = 1.0,
      tminpwl$R = 1.0,
      tminpwh$R = 1.0,
      tsetup$R$CK = 1.0,
      thold$R$CK = 0.5,
      tplh$CK$QN = 1.0,
      tphl$CK$QN = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (QN -: D)) = (tplh$CK$QN, tphl$CK$QN);
    if ( SandRandSE )
      (posedge CK *> (QN -: SI)) = (tplh$CK$QN, tphl$CK$QN);

// timing checks
    $setuphold(posedge CK, negedge R, tsetup$R$CK ,thold$R$CK , NOTIFIER);
    $width(posedge R, tminpwh$R, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 

endspecify
endmodule // SDFFRPQNX1MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFRPQNX0P5MA10TR (QN, D, SI, SE, CK, R);
output QN;
input D, SI, SE, CK, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  not     I72 (QN, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$R$QN = 1.0,
      tphl$R$QN = 1.0,
      tminpwl$R = 1.0,
      tminpwh$R = 1.0,
      tsetup$R$CK = 1.0,
      thold$R$CK = 0.5,
      tplh$CK$QN = 1.0,
      tphl$CK$QN = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (QN -: D)) = (tplh$CK$QN, tphl$CK$QN);
    if ( SandRandSE )
      (posedge CK *> (QN -: SI)) = (tplh$CK$QN, tphl$CK$QN);

// timing checks
    $setuphold(posedge CK, negedge R, tsetup$R$CK ,thold$R$CK , NOTIFIER);
    $width(posedge R, tminpwh$R, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (posedge  R *> (QN -: 1'b1)) = (tphl$R$QN); 

endspecify
endmodule // SDFFRPQNX0P5MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFRPQX4MA10TR (Q, D, SI, SE, CK, R);
output Q;
input D, SI, SE, CK, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$R$Q = 1.0,
      tphl$R$Q = 1.0,
      tminpwl$R = 1.0,
      tminpwh$R = 1.0,
      tsetup$R$CK = 1.0,
      thold$R$CK = 0.5,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK, negedge R, tsetup$R$CK ,thold$R$CK , NOTIFIER);
    $width(posedge R, tminpwh$R, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 

endspecify
endmodule // SDFFRPQX4MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFRPQX3MA10TR (Q, D, SI, SE, CK, R);
output Q;
input D, SI, SE, CK, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$R$Q = 1.0,
      tphl$R$Q = 1.0,
      tminpwl$R = 1.0,
      tminpwh$R = 1.0,
      tsetup$R$CK = 1.0,
      thold$R$CK = 0.5,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK, negedge R, tsetup$R$CK ,thold$R$CK , NOTIFIER);
    $width(posedge R, tminpwh$R, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 

endspecify
endmodule // SDFFRPQX3MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFRPQX2MA10TR (Q, D, SI, SE, CK, R);
output Q;
input D, SI, SE, CK, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$R$Q = 1.0,
      tphl$R$Q = 1.0,
      tminpwl$R = 1.0,
      tminpwh$R = 1.0,
      tsetup$R$CK = 1.0,
      thold$R$CK = 0.5,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK, negedge R, tsetup$R$CK ,thold$R$CK , NOTIFIER);
    $width(posedge R, tminpwh$R, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 

endspecify
endmodule // SDFFRPQX2MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFRPQX1MA10TR (Q, D, SI, SE, CK, R);
output Q;
input D, SI, SE, CK, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$R$Q = 1.0,
      tphl$R$Q = 1.0,
      tminpwl$R = 1.0,
      tminpwh$R = 1.0,
      tsetup$R$CK = 1.0,
      thold$R$CK = 0.5,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK, negedge R, tsetup$R$CK ,thold$R$CK , NOTIFIER);
    $width(posedge R, tminpwh$R, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 

endspecify
endmodule // SDFFRPQX1MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFRPQX0P5MA10TR (Q, D, SI, SE, CK, R);
output Q;
input D, SI, SE, CK, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$R$Q = 1.0,
      tphl$R$Q = 1.0,
      tminpwl$R = 1.0,
      tminpwh$R = 1.0,
      tsetup$R$CK = 1.0,
      thold$R$CK = 0.5,
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK, negedge R, tsetup$R$CK ,thold$R$CK , NOTIFIER);
    $width(posedge R, tminpwh$R, 0, NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 

endspecify
endmodule // SDFFRPQX0P5MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFQNX3MA10TR (QN, D, SI, SE, CK);
output QN;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  not     I72 (QN, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$CK$QN = 1.0,
      tphl$CK$QN = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (QN -: D)) = (tplh$CK$QN, tphl$CK$QN);
    if ( SandRandSE )
      (posedge CK *> (QN -: SI)) = (tplh$CK$QN, tphl$CK$QN);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // SDFFQNX3MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFQNX2MA10TR (QN, D, SI, SE, CK);
output QN;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  not     I72 (QN, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$CK$QN = 1.0,
      tphl$CK$QN = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (QN -: D)) = (tplh$CK$QN, tphl$CK$QN);
    if ( SandRandSE )
      (posedge CK *> (QN -: SI)) = (tplh$CK$QN, tphl$CK$QN);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // SDFFQNX2MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFQNX1MA10TR (QN, D, SI, SE, CK);
output QN;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  not     I72 (QN, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$CK$QN = 1.0,
      tphl$CK$QN = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (QN -: D)) = (tplh$CK$QN, tphl$CK$QN);
    if ( SandRandSE )
      (posedge CK *> (QN -: SI)) = (tplh$CK$QN, tphl$CK$QN);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // SDFFQNX1MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFQNX0P5MA10TR (QN, D, SI, SE, CK);
output QN;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  not     I72 (QN, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$CK$QN = 1.0,
      tphl$CK$QN = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (QN -: D)) = (tplh$CK$QN, tphl$CK$QN);
    if ( SandRandSE )
      (posedge CK *> (QN -: SI)) = (tplh$CK$QN, tphl$CK$QN);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // SDFFQNX0P5MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFQX4MA10TR (Q, D, SI, SE, CK);
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // SDFFQX4MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFQX3MA10TR (Q, D, SI, SE, CK);
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // SDFFQX3MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFQX2MA10TR (Q, D, SI, SE, CK);
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // SDFFQX2MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFQX1MA10TR (Q, D, SI, SE, CK);
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // SDFFQX1MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFQX0P5MA10TR (Q, D, SI, SE, CK);
output Q;
input D, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb )
      (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge D, tsetup$D$CK  ,thold$D$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // SDFFQX0P5MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFNSRPQX3MA10TR (Q, D, SI, SE, CKN, SN, R);
output Q;
input D, SI, SE, CKN, SN, R;
reg NOTIFIER;
  not   XX0 (xRN, R);
  buf   XX1 (xSN, SN);
  not     IC (clk, CKN);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$SN$Q = 1.0,
      tphl$SN$Q = 1.0,
      tplh$R$Q = 1.0,
      tphl$R$Q = 1.0,
      tminpwl$SN = 1.0,
      tminpwh$SN = 1.0,
      tminpwl$R = 1.0,
      tminpwh$R = 1.0,
      tsetup$SN$CKN = 1.0,
      thold$SN$CKN = 0.5,
      tsetup$R$CKN = 1.0,
      thold$R$CKN = 0.5,
      tplh$CKN$Q = 1.0,
      tphl$CKN$Q = 1.0,
      tsetup$D$CKN = 1.0,
      thold$D$CKN = 0.5,
      tsetup$SI$CKN = 1.0,
      thold$SI$CKN = 0.5,
      tsetup$SE$CKN = 1.0,
      thold$SE$CKN = 0.5,
      thold$R$SN = 1.0,
      thold$SN$R = 1.0,
      tminpwl$CKN = 1.0,
      tminpwh$CKN = 1.0,
      tperiod$CKN = 1.0;
 // path delays
    if (SandRandSEb)
      (negedge CKN *> (Q    +: D)) = (tplh$CKN$Q,    tphl$CKN$Q);
    if (SandRandSE)
      (negedge CKN *> (Q    +: SI)) = (tplh$CKN$Q,    tphl$CKN$Q);

// timing checks
    $setuphold(negedge CKN &&& (SandRandSEb == 1), posedge D, tsetup$D$CKN  ,thold$D$CKN  , NOTIFIER);
    $setuphold(negedge CKN &&& (SandRandSEb == 1), negedge D, tsetup$D$CKN  ,thold$D$CKN  , NOTIFIER);
    $setuphold(negedge CKN &&& (SandRandSE == 1), posedge SI, tsetup$SI$CKN ,thold$SI$CKN , NOTIFIER);
    $setuphold(negedge CKN &&& (SandRandSE == 1), negedge SI, tsetup$SI$CKN ,thold$SI$CKN , NOTIFIER);
    $setuphold(negedge CKN &&& (flag == 1), posedge SE, tsetup$SE$CKN ,thold$SE$CKN , NOTIFIER);
    $setuphold(negedge CKN &&& (flag == 1), negedge SE, tsetup$SE$CKN ,thold$SE$CKN , NOTIFIER);
    $width(negedge CKN &&& (SandR == 1), tminpwl$CKN, 0, NOTIFIER);
    $width(posedge CKN &&& (SandR == 1), tminpwh$CKN, 0, NOTIFIER);
    $period(posedge CKN &&& (SandR == 1), tperiod$CKN, NOTIFIER);
    $setuphold(negedge CKN, posedge SN, tsetup$SN$CKN ,thold$SN$CKN , NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(negedge CKN, negedge R &&& (SN == 1'b1), tsetup$R$CKN ,thold$R$CKN , NOTIFIER);
    $width(posedge R &&& (SN == 1'b1), tminpwh$R, 0, NOTIFIER);
    $hold(negedge R, negedge SN, thold$SN$R, NOTIFIER);    
    $hold(posedge SN, posedge R, thold$R$SN, NOTIFIER);    
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 

endspecify
endmodule // SDFFNSRPQX3MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFNSRPQX2MA10TR (Q, D, SI, SE, CKN, SN, R);
output Q;
input D, SI, SE, CKN, SN, R;
reg NOTIFIER;
  not   XX0 (xRN, R);
  buf   XX1 (xSN, SN);
  not     IC (clk, CKN);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$SN$Q = 1.0,
      tphl$SN$Q = 1.0,
      tplh$R$Q = 1.0,
      tphl$R$Q = 1.0,
      tminpwl$SN = 1.0,
      tminpwh$SN = 1.0,
      tminpwl$R = 1.0,
      tminpwh$R = 1.0,
      tsetup$SN$CKN = 1.0,
      thold$SN$CKN = 0.5,
      tsetup$R$CKN = 1.0,
      thold$R$CKN = 0.5,
      tplh$CKN$Q = 1.0,
      tphl$CKN$Q = 1.0,
      tsetup$D$CKN = 1.0,
      thold$D$CKN = 0.5,
      tsetup$SI$CKN = 1.0,
      thold$SI$CKN = 0.5,
      tsetup$SE$CKN = 1.0,
      thold$SE$CKN = 0.5,
      thold$R$SN = 1.0,
      thold$SN$R = 1.0,
      tminpwl$CKN = 1.0,
      tminpwh$CKN = 1.0,
      tperiod$CKN = 1.0;
 // path delays
    if (SandRandSEb)
      (negedge CKN *> (Q    +: D)) = (tplh$CKN$Q,    tphl$CKN$Q);
    if (SandRandSE)
      (negedge CKN *> (Q    +: SI)) = (tplh$CKN$Q,    tphl$CKN$Q);

// timing checks
    $setuphold(negedge CKN &&& (SandRandSEb == 1), posedge D, tsetup$D$CKN  ,thold$D$CKN  , NOTIFIER);
    $setuphold(negedge CKN &&& (SandRandSEb == 1), negedge D, tsetup$D$CKN  ,thold$D$CKN  , NOTIFIER);
    $setuphold(negedge CKN &&& (SandRandSE == 1), posedge SI, tsetup$SI$CKN ,thold$SI$CKN , NOTIFIER);
    $setuphold(negedge CKN &&& (SandRandSE == 1), negedge SI, tsetup$SI$CKN ,thold$SI$CKN , NOTIFIER);
    $setuphold(negedge CKN &&& (flag == 1), posedge SE, tsetup$SE$CKN ,thold$SE$CKN , NOTIFIER);
    $setuphold(negedge CKN &&& (flag == 1), negedge SE, tsetup$SE$CKN ,thold$SE$CKN , NOTIFIER);
    $width(negedge CKN &&& (SandR == 1), tminpwl$CKN, 0, NOTIFIER);
    $width(posedge CKN &&& (SandR == 1), tminpwh$CKN, 0, NOTIFIER);
    $period(posedge CKN &&& (SandR == 1), tperiod$CKN, NOTIFIER);
    $setuphold(negedge CKN, posedge SN, tsetup$SN$CKN ,thold$SN$CKN , NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(negedge CKN, negedge R &&& (SN == 1'b1), tsetup$R$CKN ,thold$R$CKN , NOTIFIER);
    $width(posedge R &&& (SN == 1'b1), tminpwh$R, 0, NOTIFIER);
    $hold(negedge R, negedge SN, thold$SN$R, NOTIFIER);    
    $hold(posedge SN, posedge R, thold$R$SN, NOTIFIER);    
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 

endspecify
endmodule // SDFFNSRPQX2MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFNSRPQX1MA10TR (Q, D, SI, SE, CKN, SN, R);
output Q;
input D, SI, SE, CKN, SN, R;
reg NOTIFIER;
  not   XX0 (xRN, R);
  buf   XX1 (xSN, SN);
  not     IC (clk, CKN);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$SN$Q = 1.0,
      tphl$SN$Q = 1.0,
      tplh$R$Q = 1.0,
      tphl$R$Q = 1.0,
      tminpwl$SN = 1.0,
      tminpwh$SN = 1.0,
      tminpwl$R = 1.0,
      tminpwh$R = 1.0,
      tsetup$SN$CKN = 1.0,
      thold$SN$CKN = 0.5,
      tsetup$R$CKN = 1.0,
      thold$R$CKN = 0.5,
      tplh$CKN$Q = 1.0,
      tphl$CKN$Q = 1.0,
      tsetup$D$CKN = 1.0,
      thold$D$CKN = 0.5,
      tsetup$SI$CKN = 1.0,
      thold$SI$CKN = 0.5,
      tsetup$SE$CKN = 1.0,
      thold$SE$CKN = 0.5,
      thold$R$SN = 1.0,
      thold$SN$R = 1.0,
      tminpwl$CKN = 1.0,
      tminpwh$CKN = 1.0,
      tperiod$CKN = 1.0;
 // path delays
    if (SandRandSEb)
      (negedge CKN *> (Q    +: D)) = (tplh$CKN$Q,    tphl$CKN$Q);
    if (SandRandSE)
      (negedge CKN *> (Q    +: SI)) = (tplh$CKN$Q,    tphl$CKN$Q);

// timing checks
    $setuphold(negedge CKN &&& (SandRandSEb == 1), posedge D, tsetup$D$CKN  ,thold$D$CKN  , NOTIFIER);
    $setuphold(negedge CKN &&& (SandRandSEb == 1), negedge D, tsetup$D$CKN  ,thold$D$CKN  , NOTIFIER);
    $setuphold(negedge CKN &&& (SandRandSE == 1), posedge SI, tsetup$SI$CKN ,thold$SI$CKN , NOTIFIER);
    $setuphold(negedge CKN &&& (SandRandSE == 1), negedge SI, tsetup$SI$CKN ,thold$SI$CKN , NOTIFIER);
    $setuphold(negedge CKN &&& (flag == 1), posedge SE, tsetup$SE$CKN ,thold$SE$CKN , NOTIFIER);
    $setuphold(negedge CKN &&& (flag == 1), negedge SE, tsetup$SE$CKN ,thold$SE$CKN , NOTIFIER);
    $width(negedge CKN &&& (SandR == 1), tminpwl$CKN, 0, NOTIFIER);
    $width(posedge CKN &&& (SandR == 1), tminpwh$CKN, 0, NOTIFIER);
    $period(posedge CKN &&& (SandR == 1), tperiod$CKN, NOTIFIER);
    $setuphold(negedge CKN, posedge SN, tsetup$SN$CKN ,thold$SN$CKN , NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $setuphold(negedge CKN, negedge R &&& (SN == 1'b1), tsetup$R$CKN ,thold$R$CKN , NOTIFIER);
    $width(posedge R &&& (SN == 1'b1), tminpwh$R, 0, NOTIFIER);
    $hold(negedge R, negedge SN, thold$SN$R, NOTIFIER);    
    $hold(posedge SN, posedge R, thold$R$SN, NOTIFIER);    
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 && SN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 && R == 1'b0)
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 

endspecify
endmodule // SDFFNSRPQX1MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFNSQX3MA10TR (Q, D, SI, SE, CKN, SN);
output Q;
input D, SI, SE, CKN, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  not     IC (clk, CKN);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$SN$Q = 1.0,
      tphl$SN$Q = 1.0,
      tminpwl$SN = 1.0,
      tminpwh$SN = 1.0,
      tsetup$SN$CKN = 1.0,
      thold$SN$CKN = 0.5,
      tplh$CKN$Q = 1.0,
      tphl$CKN$Q = 1.0,
      tsetup$D$CKN = 1.0,
      thold$D$CKN = 0.5,
      tsetup$SI$CKN = 1.0,
      thold$SI$CKN = 0.5,
      tsetup$SE$CKN = 1.0,
      thold$SE$CKN = 0.5,
      tminpwl$CKN = 1.0,
      tminpwh$CKN = 1.0,
      tperiod$CKN = 1.0;
 // path delays
    if (SandRandSEb)
      (negedge CKN *> (Q    +: D)) = (tplh$CKN$Q,    tphl$CKN$Q);
    if (SandRandSE)
      (negedge CKN *> (Q    +: SI)) = (tplh$CKN$Q,    tphl$CKN$Q);

// timing checks
    $setuphold(negedge CKN &&& (SandRandSEb == 1), posedge D, tsetup$D$CKN  ,thold$D$CKN  , NOTIFIER);
    $setuphold(negedge CKN &&& (SandRandSEb == 1), negedge D, tsetup$D$CKN  ,thold$D$CKN  , NOTIFIER);
    $setuphold(negedge CKN &&& (SandRandSE == 1), posedge SI, tsetup$SI$CKN ,thold$SI$CKN , NOTIFIER);
    $setuphold(negedge CKN &&& (SandRandSE == 1), negedge SI, tsetup$SI$CKN ,thold$SI$CKN , NOTIFIER);
    $setuphold(negedge CKN &&& (flag == 1), posedge SE, tsetup$SE$CKN ,thold$SE$CKN , NOTIFIER);
    $setuphold(negedge CKN &&& (flag == 1), negedge SE, tsetup$SE$CKN ,thold$SE$CKN , NOTIFIER);
    $width(negedge CKN &&& (SandR == 1), tminpwl$CKN, 0, NOTIFIER);
    $width(posedge CKN &&& (SandR == 1), tminpwh$CKN, 0, NOTIFIER);
    $period(posedge CKN &&& (SandR == 1), tperiod$CKN, NOTIFIER);
    $setuphold(negedge CKN, posedge SN, tsetup$SN$CKN ,thold$SN$CKN , NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 

endspecify
endmodule // SDFFNSQX3MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFNSQX2MA10TR (Q, D, SI, SE, CKN, SN);
output Q;
input D, SI, SE, CKN, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  not     IC (clk, CKN);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$SN$Q = 1.0,
      tphl$SN$Q = 1.0,
      tminpwl$SN = 1.0,
      tminpwh$SN = 1.0,
      tsetup$SN$CKN = 1.0,
      thold$SN$CKN = 0.5,
      tplh$CKN$Q = 1.0,
      tphl$CKN$Q = 1.0,
      tsetup$D$CKN = 1.0,
      thold$D$CKN = 0.5,
      tsetup$SI$CKN = 1.0,
      thold$SI$CKN = 0.5,
      tsetup$SE$CKN = 1.0,
      thold$SE$CKN = 0.5,
      tminpwl$CKN = 1.0,
      tminpwh$CKN = 1.0,
      tperiod$CKN = 1.0;
 // path delays
    if (SandRandSEb)
      (negedge CKN *> (Q    +: D)) = (tplh$CKN$Q,    tphl$CKN$Q);
    if (SandRandSE)
      (negedge CKN *> (Q    +: SI)) = (tplh$CKN$Q,    tphl$CKN$Q);

// timing checks
    $setuphold(negedge CKN &&& (SandRandSEb == 1), posedge D, tsetup$D$CKN  ,thold$D$CKN  , NOTIFIER);
    $setuphold(negedge CKN &&& (SandRandSEb == 1), negedge D, tsetup$D$CKN  ,thold$D$CKN  , NOTIFIER);
    $setuphold(negedge CKN &&& (SandRandSE == 1), posedge SI, tsetup$SI$CKN ,thold$SI$CKN , NOTIFIER);
    $setuphold(negedge CKN &&& (SandRandSE == 1), negedge SI, tsetup$SI$CKN ,thold$SI$CKN , NOTIFIER);
    $setuphold(negedge CKN &&& (flag == 1), posedge SE, tsetup$SE$CKN ,thold$SE$CKN , NOTIFIER);
    $setuphold(negedge CKN &&& (flag == 1), negedge SE, tsetup$SE$CKN ,thold$SE$CKN , NOTIFIER);
    $width(negedge CKN &&& (SandR == 1), tminpwl$CKN, 0, NOTIFIER);
    $width(posedge CKN &&& (SandR == 1), tminpwh$CKN, 0, NOTIFIER);
    $period(posedge CKN &&& (SandR == 1), tperiod$CKN, NOTIFIER);
    $setuphold(negedge CKN, posedge SN, tsetup$SN$CKN ,thold$SN$CKN , NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 

endspecify
endmodule // SDFFNSQX2MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFNSQX1MA10TR (Q, D, SI, SE, CKN, SN);
output Q;
input D, SI, SE, CKN, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

  buf   XX0 (xSN, SN);
  not     IC (clk, CKN);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$SN$Q = 1.0,
      tphl$SN$Q = 1.0,
      tminpwl$SN = 1.0,
      tminpwh$SN = 1.0,
      tsetup$SN$CKN = 1.0,
      thold$SN$CKN = 0.5,
      tplh$CKN$Q = 1.0,
      tphl$CKN$Q = 1.0,
      tsetup$D$CKN = 1.0,
      thold$D$CKN = 0.5,
      tsetup$SI$CKN = 1.0,
      thold$SI$CKN = 0.5,
      tsetup$SE$CKN = 1.0,
      thold$SE$CKN = 0.5,
      tminpwl$CKN = 1.0,
      tminpwh$CKN = 1.0,
      tperiod$CKN = 1.0;
 // path delays
    if (SandRandSEb)
      (negedge CKN *> (Q    +: D)) = (tplh$CKN$Q,    tphl$CKN$Q);
    if (SandRandSE)
      (negedge CKN *> (Q    +: SI)) = (tplh$CKN$Q,    tphl$CKN$Q);

// timing checks
    $setuphold(negedge CKN &&& (SandRandSEb == 1), posedge D, tsetup$D$CKN  ,thold$D$CKN  , NOTIFIER);
    $setuphold(negedge CKN &&& (SandRandSEb == 1), negedge D, tsetup$D$CKN  ,thold$D$CKN  , NOTIFIER);
    $setuphold(negedge CKN &&& (SandRandSE == 1), posedge SI, tsetup$SI$CKN ,thold$SI$CKN , NOTIFIER);
    $setuphold(negedge CKN &&& (SandRandSE == 1), negedge SI, tsetup$SI$CKN ,thold$SI$CKN , NOTIFIER);
    $setuphold(negedge CKN &&& (flag == 1), posedge SE, tsetup$SE$CKN ,thold$SE$CKN , NOTIFIER);
    $setuphold(negedge CKN &&& (flag == 1), negedge SE, tsetup$SE$CKN ,thold$SE$CKN , NOTIFIER);
    $width(negedge CKN &&& (SandR == 1), tminpwl$CKN, 0, NOTIFIER);
    $width(posedge CKN &&& (SandR == 1), tminpwh$CKN, 0, NOTIFIER);
    $period(posedge CKN &&& (SandR == 1), tperiod$CKN, NOTIFIER);
    $setuphold(negedge CKN, posedge SN, tsetup$SN$CKN ,thold$SN$CKN , NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 )
       (negedge  SN *> (Q +: 1'b0)) = (tplh$SN$Q); 

endspecify
endmodule // SDFFNSQX1MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFNRPQX3MA10TR (Q, D, SI, SE, CKN, R);
output Q;
input D, SI, SE, CKN, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  not     IC (clk, CKN);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$R$Q = 1.0,
      tphl$R$Q = 1.0,
      tminpwl$R = 1.0,
      tminpwh$R = 1.0,
      tsetup$R$CKN = 1.0,
      thold$R$CKN = 0.5,
      tplh$CKN$Q = 1.0,
      tphl$CKN$Q = 1.0,
      tsetup$D$CKN = 1.0,
      thold$D$CKN = 0.5,
      tsetup$SI$CKN = 1.0,
      thold$SI$CKN = 0.5,
      tsetup$SE$CKN = 1.0,
      thold$SE$CKN = 0.5,
      tminpwl$CKN = 1.0,
      tminpwh$CKN = 1.0,
      tperiod$CKN = 1.0;
 // path delays
    if (SandRandSEb)
      (negedge CKN *> (Q    +: D)) = (tplh$CKN$Q,    tphl$CKN$Q);
    if (SandRandSE)
      (negedge CKN *> (Q    +: SI)) = (tplh$CKN$Q,    tphl$CKN$Q);

// timing checks
    $setuphold(negedge CKN &&& (SandRandSEb == 1), posedge D, tsetup$D$CKN  ,thold$D$CKN  , NOTIFIER);
    $setuphold(negedge CKN &&& (SandRandSEb == 1), negedge D, tsetup$D$CKN  ,thold$D$CKN  , NOTIFIER);
    $setuphold(negedge CKN &&& (SandRandSE == 1), posedge SI, tsetup$SI$CKN ,thold$SI$CKN , NOTIFIER);
    $setuphold(negedge CKN &&& (SandRandSE == 1), negedge SI, tsetup$SI$CKN ,thold$SI$CKN , NOTIFIER);
    $setuphold(negedge CKN &&& (flag == 1), posedge SE, tsetup$SE$CKN ,thold$SE$CKN , NOTIFIER);
    $setuphold(negedge CKN &&& (flag == 1), negedge SE, tsetup$SE$CKN ,thold$SE$CKN , NOTIFIER);
    $setuphold(negedge CKN, negedge R, tsetup$R$CKN ,thold$R$CKN , NOTIFIER);
    $width(posedge R, tminpwh$R, 0, NOTIFIER);
    $width(negedge CKN &&& (SandR == 1), tminpwl$CKN, 0, NOTIFIER);
    $width(posedge CKN &&& (SandR == 1), tminpwh$CKN, 0, NOTIFIER);
    $period(posedge CKN &&& (SandR == 1), tperiod$CKN, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 

endspecify
endmodule // SDFFNRPQX3MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFNRPQX2MA10TR (Q, D, SI, SE, CKN, R);
output Q;
input D, SI, SE, CKN, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  not     IC (clk, CKN);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$R$Q = 1.0,
      tphl$R$Q = 1.0,
      tminpwl$R = 1.0,
      tminpwh$R = 1.0,
      tsetup$R$CKN = 1.0,
      thold$R$CKN = 0.5,
      tplh$CKN$Q = 1.0,
      tphl$CKN$Q = 1.0,
      tsetup$D$CKN = 1.0,
      thold$D$CKN = 0.5,
      tsetup$SI$CKN = 1.0,
      thold$SI$CKN = 0.5,
      tsetup$SE$CKN = 1.0,
      thold$SE$CKN = 0.5,
      tminpwl$CKN = 1.0,
      tminpwh$CKN = 1.0,
      tperiod$CKN = 1.0;
 // path delays
    if (SandRandSEb)
      (negedge CKN *> (Q    +: D)) = (tplh$CKN$Q,    tphl$CKN$Q);
    if (SandRandSE)
      (negedge CKN *> (Q    +: SI)) = (tplh$CKN$Q,    tphl$CKN$Q);

// timing checks
    $setuphold(negedge CKN &&& (SandRandSEb == 1), posedge D, tsetup$D$CKN  ,thold$D$CKN  , NOTIFIER);
    $setuphold(negedge CKN &&& (SandRandSEb == 1), negedge D, tsetup$D$CKN  ,thold$D$CKN  , NOTIFIER);
    $setuphold(negedge CKN &&& (SandRandSE == 1), posedge SI, tsetup$SI$CKN ,thold$SI$CKN , NOTIFIER);
    $setuphold(negedge CKN &&& (SandRandSE == 1), negedge SI, tsetup$SI$CKN ,thold$SI$CKN , NOTIFIER);
    $setuphold(negedge CKN &&& (flag == 1), posedge SE, tsetup$SE$CKN ,thold$SE$CKN , NOTIFIER);
    $setuphold(negedge CKN &&& (flag == 1), negedge SE, tsetup$SE$CKN ,thold$SE$CKN , NOTIFIER);
    $setuphold(negedge CKN, negedge R, tsetup$R$CKN ,thold$R$CKN , NOTIFIER);
    $width(posedge R, tminpwh$R, 0, NOTIFIER);
    $width(negedge CKN &&& (SandR == 1), tminpwl$CKN, 0, NOTIFIER);
    $width(posedge CKN &&& (SandR == 1), tminpwh$CKN, 0, NOTIFIER);
    $period(posedge CKN &&& (SandR == 1), tperiod$CKN, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 

endspecify
endmodule // SDFFNRPQX2MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFNRPQX1MA10TR (Q, D, SI, SE, CKN, R);
output Q;
input D, SI, SE, CKN, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

  not   XX0 (xRN, R); 
  not     IC (clk, CKN);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$R$Q = 1.0,
      tphl$R$Q = 1.0,
      tminpwl$R = 1.0,
      tminpwh$R = 1.0,
      tsetup$R$CKN = 1.0,
      thold$R$CKN = 0.5,
      tplh$CKN$Q = 1.0,
      tphl$CKN$Q = 1.0,
      tsetup$D$CKN = 1.0,
      thold$D$CKN = 0.5,
      tsetup$SI$CKN = 1.0,
      thold$SI$CKN = 0.5,
      tsetup$SE$CKN = 1.0,
      thold$SE$CKN = 0.5,
      tminpwl$CKN = 1.0,
      tminpwh$CKN = 1.0,
      tperiod$CKN = 1.0;
 // path delays
    if (SandRandSEb)
      (negedge CKN *> (Q    +: D)) = (tplh$CKN$Q,    tphl$CKN$Q);
    if (SandRandSE)
      (negedge CKN *> (Q    +: SI)) = (tplh$CKN$Q,    tphl$CKN$Q);

// timing checks
    $setuphold(negedge CKN &&& (SandRandSEb == 1), posedge D, tsetup$D$CKN  ,thold$D$CKN  , NOTIFIER);
    $setuphold(negedge CKN &&& (SandRandSEb == 1), negedge D, tsetup$D$CKN  ,thold$D$CKN  , NOTIFIER);
    $setuphold(negedge CKN &&& (SandRandSE == 1), posedge SI, tsetup$SI$CKN ,thold$SI$CKN , NOTIFIER);
    $setuphold(negedge CKN &&& (SandRandSE == 1), negedge SI, tsetup$SI$CKN ,thold$SI$CKN , NOTIFIER);
    $setuphold(negedge CKN &&& (flag == 1), posedge SE, tsetup$SE$CKN ,thold$SE$CKN , NOTIFIER);
    $setuphold(negedge CKN &&& (flag == 1), negedge SE, tsetup$SE$CKN ,thold$SE$CKN , NOTIFIER);
    $setuphold(negedge CKN, negedge R, tsetup$R$CKN ,thold$R$CKN , NOTIFIER);
    $width(posedge R, tminpwh$R, 0, NOTIFIER);
    $width(negedge CKN &&& (SandR == 1), tminpwl$CKN, 0, NOTIFIER);
    $width(posedge CKN &&& (SandR == 1), tminpwh$CKN, 0, NOTIFIER);
    $period(posedge CKN &&& (SandR == 1), tperiod$CKN, NOTIFIER);
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b0 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b0 && CKN == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b0 && D == 1'b1 && CKN == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b0 && CKN == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 
    if (SI == 1'b1 && SE == 1'b1 && D == 1'b1 && CKN == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = (tphl$R$Q); 

endspecify
endmodule // SDFFNRPQX1MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFNQX3MA10TR (Q, D, SI, SE, CKN);
output Q;
input D, SI, SE, CKN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  not     IC (clk, CKN);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$CKN$Q = 1.0,
      tphl$CKN$Q = 1.0,
      tsetup$D$CKN = 1.0,
      thold$D$CKN = 0.5,
      tsetup$SI$CKN = 1.0,
      thold$SI$CKN = 0.5,
      tsetup$SE$CKN = 1.0,
      thold$SE$CKN = 0.5,
      tminpwl$CKN = 1.0,
      tminpwh$CKN = 1.0,
      tperiod$CKN = 1.0;
 // path delays
    if (SandRandSEb)
      (negedge CKN *> (Q    +: D)) = (tplh$CKN$Q,    tphl$CKN$Q);
    if (SandRandSE)
      (negedge CKN *> (Q    +: SI)) = (tplh$CKN$Q,    tphl$CKN$Q);

// timing checks
    $setuphold(negedge CKN &&& (SandRandSEb == 1), posedge D, tsetup$D$CKN  ,thold$D$CKN  , NOTIFIER);
    $setuphold(negedge CKN &&& (SandRandSEb == 1), negedge D, tsetup$D$CKN  ,thold$D$CKN  , NOTIFIER);
    $setuphold(negedge CKN &&& (SandRandSE == 1), posedge SI, tsetup$SI$CKN ,thold$SI$CKN , NOTIFIER);
    $setuphold(negedge CKN &&& (SandRandSE == 1), negedge SI, tsetup$SI$CKN ,thold$SI$CKN , NOTIFIER);
    $setuphold(negedge CKN &&& (flag == 1), posedge SE, tsetup$SE$CKN ,thold$SE$CKN , NOTIFIER);
    $setuphold(negedge CKN &&& (flag == 1), negedge SE, tsetup$SE$CKN ,thold$SE$CKN , NOTIFIER);
    $width(negedge CKN &&& (SandR == 1), tminpwl$CKN, 0, NOTIFIER);
    $width(posedge CKN &&& (SandR == 1), tminpwh$CKN, 0, NOTIFIER);
    $period(posedge CKN &&& (SandR == 1), tperiod$CKN, NOTIFIER);

endspecify
endmodule // SDFFNQX3MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFNQX2MA10TR (Q, D, SI, SE, CKN);
output Q;
input D, SI, SE, CKN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  not     IC (clk, CKN);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$CKN$Q = 1.0,
      tphl$CKN$Q = 1.0,
      tsetup$D$CKN = 1.0,
      thold$D$CKN = 0.5,
      tsetup$SI$CKN = 1.0,
      thold$SI$CKN = 0.5,
      tsetup$SE$CKN = 1.0,
      thold$SE$CKN = 0.5,
      tminpwl$CKN = 1.0,
      tminpwh$CKN = 1.0,
      tperiod$CKN = 1.0;
 // path delays
    if (SandRandSEb)
      (negedge CKN *> (Q    +: D)) = (tplh$CKN$Q,    tphl$CKN$Q);
    if (SandRandSE)
      (negedge CKN *> (Q    +: SI)) = (tplh$CKN$Q,    tphl$CKN$Q);

// timing checks
    $setuphold(negedge CKN &&& (SandRandSEb == 1), posedge D, tsetup$D$CKN  ,thold$D$CKN  , NOTIFIER);
    $setuphold(negedge CKN &&& (SandRandSEb == 1), negedge D, tsetup$D$CKN  ,thold$D$CKN  , NOTIFIER);
    $setuphold(negedge CKN &&& (SandRandSE == 1), posedge SI, tsetup$SI$CKN ,thold$SI$CKN , NOTIFIER);
    $setuphold(negedge CKN &&& (SandRandSE == 1), negedge SI, tsetup$SI$CKN ,thold$SI$CKN , NOTIFIER);
    $setuphold(negedge CKN &&& (flag == 1), posedge SE, tsetup$SE$CKN ,thold$SE$CKN , NOTIFIER);
    $setuphold(negedge CKN &&& (flag == 1), negedge SE, tsetup$SE$CKN ,thold$SE$CKN , NOTIFIER);
    $width(negedge CKN &&& (SandR == 1), tminpwl$CKN, 0, NOTIFIER);
    $width(posedge CKN &&& (SandR == 1), tminpwh$CKN, 0, NOTIFIER);
    $period(posedge CKN &&& (SandR == 1), tperiod$CKN, NOTIFIER);

endspecify
endmodule // SDFFNQX2MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module SDFFNQX1MA10TR (Q, D, SI, SE, CKN);
output Q;
input D, SI, SE, CKN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  not     IC (clk, CKN);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I1 (n1, D, SI, SE);
  buf     I2 (Q, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  xor     I8 (DxorSD, D, SI);
  and     I9 (flag, DxorSD, SandR);
  specify
    specparam 
      tplh$CKN$Q = 1.0,
      tphl$CKN$Q = 1.0,
      tsetup$D$CKN = 1.0,
      thold$D$CKN = 0.5,
      tsetup$SI$CKN = 1.0,
      thold$SI$CKN = 0.5,
      tsetup$SE$CKN = 1.0,
      thold$SE$CKN = 0.5,
      tminpwl$CKN = 1.0,
      tminpwh$CKN = 1.0,
      tperiod$CKN = 1.0;
 // path delays
    if (SandRandSEb)
      (negedge CKN *> (Q    +: D)) = (tplh$CKN$Q,    tphl$CKN$Q);
    if (SandRandSE)
      (negedge CKN *> (Q    +: SI)) = (tplh$CKN$Q,    tphl$CKN$Q);

// timing checks
    $setuphold(negedge CKN &&& (SandRandSEb == 1), posedge D, tsetup$D$CKN  ,thold$D$CKN  , NOTIFIER);
    $setuphold(negedge CKN &&& (SandRandSEb == 1), negedge D, tsetup$D$CKN  ,thold$D$CKN  , NOTIFIER);
    $setuphold(negedge CKN &&& (SandRandSE == 1), posedge SI, tsetup$SI$CKN ,thold$SI$CKN , NOTIFIER);
    $setuphold(negedge CKN &&& (SandRandSE == 1), negedge SI, tsetup$SI$CKN ,thold$SI$CKN , NOTIFIER);
    $setuphold(negedge CKN &&& (flag == 1), posedge SE, tsetup$SE$CKN ,thold$SE$CKN , NOTIFIER);
    $setuphold(negedge CKN &&& (flag == 1), negedge SE, tsetup$SE$CKN ,thold$SE$CKN , NOTIFIER);
    $width(negedge CKN &&& (SandR == 1), tminpwl$CKN, 0, NOTIFIER);
    $width(posedge CKN &&& (SandR == 1), tminpwh$CKN, 0, NOTIFIER);
    $period(posedge CKN &&& (SandR == 1), tperiod$CKN, NOTIFIER);

endspecify
endmodule // SDFFNQX1MA10TR
`endcelldefine
	

//$Id: rf.genpp,v 1.11 2006/05/18 09:44:11 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module RF2R2WSX2MA10TR (RBL1, RBL2, WBL1, WWL1, WBL2, WWL2, RWL1, RWL2);
output RBL1, RBL2;
input WBL1, WWL1, WBL2, WWL2, RWL1, RWL2;
reg NOTIFIER;

   or  I0 (ck, WWL1, WWL2);
   not I1 (ckn, ck);
   udp_wao I2 (wr, WBL1, WBL2, WWL1, WWL2);
   udp_tlatrf I3 (n0, wr, ck, ckn, NOTIFIER);
   not I4 (n1, n0);
   notif1 I5 (RBL1, n1, RWL1);
   notif1 I6 (RBL2, n1, RWL2);

  specify
    // delay parameters
    specparam
      tplh$WBL1$RBL1 = 1.0,
      tphl$WBL1$RBL1 = 1.0,
      tpxh$WBL1$RBL1 = 1.0,
      tphx$WBL1$RBL1 = 1.0,
      tplx$WBL1$RBL1 = 1.0,
      tpxl$WBL1$RBL1 = 1.0,
      tplh$WWL1$RBL1 = 1.0,
      tphl$WWL1$RBL1 = 1.0,
      tpxh$WWL1$RBL1 = 1.0,
      tphx$WWL1$RBL1 = 1.0,
      tplx$WWL1$RBL1 = 1.0,
      tpxl$WWL1$RBL1 = 1.0,
      tplh$WBL2$RBL1 = 1.0,
      tphl$WBL2$RBL1 = 1.0,
      tpxh$WBL2$RBL1 = 1.0,
      tphx$WBL2$RBL1 = 1.0,
      tplx$WBL2$RBL1 = 1.0,
      tpxl$WBL2$RBL1 = 1.0,
      tplh$WWL2$RBL1 = 1.0,
      tphl$WWL2$RBL1 = 1.0,
      tpxh$WWL2$RBL1 = 1.0,
      tphx$WWL2$RBL1 = 1.0,
      tplx$WWL2$RBL1 = 1.0,
      tpxl$WWL2$RBL1 = 1.0,
      tplh$RWL1$RBL1 = 1.0,
      tphl$RWL1$RBL1 = 1.0,
      tpxh$RWL1$RBL1 = 1.0,
      tphx$RWL1$RBL1 = 1.0,
      tplx$RWL1$RBL1 = 1.0,
      tpxl$RWL1$RBL1 = 1.0,
      tplh$RWL2$RBL1 = 1.0,
      tphl$RWL2$RBL1 = 1.0,
      tpxh$RWL2$RBL1 = 1.0,
      tphx$RWL2$RBL1 = 1.0,
      tplx$RWL2$RBL1 = 1.0,
      tpxl$RWL2$RBL1 = 1.0,
      tplh$WBL1$RBL2 = 1.0,
      tphl$WBL1$RBL2 = 1.0,
      tpxh$WBL1$RBL2 = 1.0,
      tphx$WBL1$RBL2 = 1.0,
      tplx$WBL1$RBL2 = 1.0,
      tpxl$WBL1$RBL2 = 1.0,
      tplh$WWL1$RBL2 = 1.0,
      tphl$WWL1$RBL2 = 1.0,
      tpxh$WWL1$RBL2 = 1.0,
      tphx$WWL1$RBL2 = 1.0,
      tplx$WWL1$RBL2 = 1.0,
      tpxl$WWL1$RBL2 = 1.0,
      tplh$WBL2$RBL2 = 1.0,
      tphl$WBL2$RBL2 = 1.0,
      tpxh$WBL2$RBL2 = 1.0,
      tphx$WBL2$RBL2 = 1.0,
      tplx$WBL2$RBL2 = 1.0,
      tpxl$WBL2$RBL2 = 1.0,
      tplh$WWL2$RBL2 = 1.0,
      tphl$WWL2$RBL2 = 1.0,
      tpxh$WWL2$RBL2 = 1.0,
      tphx$WWL2$RBL2 = 1.0,
      tplx$WWL2$RBL2 = 1.0,
      tpxl$WWL2$RBL2 = 1.0,
      tplh$RWL1$RBL2 = 1.0,
      tphl$RWL1$RBL2 = 1.0,
      tpxh$RWL1$RBL2 = 1.0,
      tphx$RWL1$RBL2 = 1.0,
      tplx$RWL1$RBL2 = 1.0,
      tpxl$RWL1$RBL2 = 1.0,
      tplh$RWL2$RBL2 = 1.0,
      tphl$RWL2$RBL2 = 1.0,
      tpxh$RWL2$RBL2 = 1.0,
      tphx$RWL2$RBL2 = 1.0,
      tplx$RWL2$RBL2 = 1.0,
      tpxl$RWL2$RBL2 = 1.0,
    tminpwh$WWL1    = 1.0,
    tperiod$WWL1    = 1.0,
    tminpwh$WWL2    = 1.0,
    tperiod$WWL2    = 1.0,
    tsetup$WWL1$WBL1 = 1.0,
    thold$WWL1$WBL1  = 0.5,
    tsetup$WWL2$WBL2 = 1.0,
    thold$WWL2$WBL2  = 0.5;

      // path delays
 
      // timing checks
      $setuphold(negedge WWL1, posedge WBL1, tsetup$WWL1$WBL1, thold$WWL1$WBL1, NOTIFIER);
      $setuphold(negedge WWL1, negedge WBL1, tsetup$WWL1$WBL1, thold$WWL1$WBL1, NOTIFIER);
      $setuphold(negedge WWL2, posedge WBL2, tsetup$WWL2$WBL2, thold$WWL2$WBL2, NOTIFIER);
      $setuphold(negedge WWL2, negedge WBL2, tsetup$WWL2$WBL2, thold$WWL2$WBL2, NOTIFIER);
      $width(posedge WWL1, tminpwh$WWL1, 0, NOTIFIER);
      $period(posedge WWL1, tperiod$WWL1, NOTIFIER);
      $width(posedge WWL2, tminpwh$WWL2, 0, NOTIFIER);
      $period(posedge WWL2, tperiod$WWL2, NOTIFIER);
    if (WWL1==1'b0 && WWL2==1'b0 && RWL2==1'b0 )
       (RWL1 *> RBL1) = (tplh$RWL1$RBL1, tphl$RWL1$RBL1, tpxh$RWL1$RBL1, tphx$RWL1$RBL1, tplx$RWL1$RBL1, tpxl$RWL1$RBL1);
    if (WWL1==1'b0 && WWL2==1'b0 && RWL1==1'b0 )
       (RWL2 *> RBL2) = (tplh$RWL2$RBL2, tphl$RWL2$RBL2, tpxh$RWL2$RBL2, tphx$RWL2$RBL2, tplx$RWL2$RBL2, tpxl$RWL2$RBL2);
    if (WWL1==1'b0 && WWL2==1'b0 && RWL2==1'b1 )
       (RWL1 *> RBL1) = (tplh$RWL1$RBL1, tphl$RWL1$RBL1, tpxh$RWL1$RBL1, tphx$RWL1$RBL1, tplx$RWL1$RBL1, tpxl$RWL1$RBL1);
    if (WWL1==1'b0 && WWL2==1'b0 && RWL1==1'b1 )
       (RWL2 *> RBL2) = (tplh$RWL2$RBL2, tphl$RWL2$RBL2, tpxh$RWL2$RBL2, tphx$RWL2$RBL2, tplx$RWL2$RBL2, tpxl$RWL2$RBL2);
    if (WWL1==1'b0 && WWL2==1'b1 && RWL2==1'b0 )
       (RWL1 *> RBL1) = (tplh$RWL1$RBL1, tphl$RWL1$RBL1, tpxh$RWL1$RBL1, tphx$RWL1$RBL1, tplx$RWL1$RBL1, tpxl$RWL1$RBL1);
    if (WWL1==1'b0 && WWL2==1'b1 && RWL1==1'b0 )
       (RWL2 *> RBL2) = (tplh$RWL2$RBL2, tphl$RWL2$RBL2, tpxh$RWL2$RBL2, tphx$RWL2$RBL2, tplx$RWL2$RBL2, tpxl$RWL2$RBL2);
    if (WWL1==1'b0 && WWL2==1'b1 && RWL2==1'b1 )
       (RWL1 *> RBL1) = (tplh$RWL1$RBL1, tphl$RWL1$RBL1, tpxh$RWL1$RBL1, tphx$RWL1$RBL1, tplx$RWL1$RBL1, tpxl$RWL1$RBL1);
    if (WWL1==1'b0 && WWL2==1'b1 && RWL1==1'b1 )
       (RWL2 *> RBL2) = (tplh$RWL2$RBL2, tphl$RWL2$RBL2, tpxh$RWL2$RBL2, tphx$RWL2$RBL2, tplx$RWL2$RBL2, tpxl$RWL2$RBL2);
    if (WWL1==1'b1 && WWL2==1'b0 && RWL2==1'b0 )
       (RWL1 *> RBL1) = (tplh$RWL1$RBL1, tphl$RWL1$RBL1, tpxh$RWL1$RBL1, tphx$RWL1$RBL1, tplx$RWL1$RBL1, tpxl$RWL1$RBL1);
    if (WWL1==1'b1 && WWL2==1'b0 && RWL1==1'b0 )
       (RWL2 *> RBL2) = (tplh$RWL2$RBL2, tphl$RWL2$RBL2, tpxh$RWL2$RBL2, tphx$RWL2$RBL2, tplx$RWL2$RBL2, tpxl$RWL2$RBL2);
    if (WWL1==1'b1 && WWL2==1'b0 && RWL2==1'b1 )
       (RWL1 *> RBL1) = (tplh$RWL1$RBL1, tphl$RWL1$RBL1, tpxh$RWL1$RBL1, tphx$RWL1$RBL1, tplx$RWL1$RBL1, tpxl$RWL1$RBL1);
    if (WWL1==1'b1 && WWL2==1'b0 && RWL1==1'b1 )
       (RWL2 *> RBL2) = (tplh$RWL2$RBL2, tphl$RWL2$RBL2, tpxh$RWL2$RBL2, tphx$RWL2$RBL2, tplx$RWL2$RBL2, tpxl$RWL2$RBL2);
    if (WWL1==1'b1 && WWL2==1'b1 && RWL2==1'b0 )
       (RWL1 *> RBL1) = (tplh$RWL1$RBL1, tphl$RWL1$RBL1, tpxh$RWL1$RBL1, tphx$RWL1$RBL1, tplx$RWL1$RBL1, tpxl$RWL1$RBL1);
    if (WWL1==1'b1 && WWL2==1'b1 && RWL1==1'b0 )
       (RWL2 *> RBL2) = (tplh$RWL2$RBL2, tphl$RWL2$RBL2, tpxh$RWL2$RBL2, tphx$RWL2$RBL2, tplx$RWL2$RBL2, tpxl$RWL2$RBL2);
    if (WWL1==1'b1 && WWL2==1'b1 && RWL2==1'b1 )
       (RWL1 *> RBL1) = (tplh$RWL1$RBL1, tphl$RWL1$RBL1, tpxh$RWL1$RBL1, tphx$RWL1$RBL1, tplx$RWL1$RBL1, tpxl$RWL1$RBL1);
    if (WWL1==1'b1 && WWL2==1'b1 && RWL1==1'b1 )
       (RWL2 *> RBL2) = (tplh$RWL2$RBL2, tphl$RWL2$RBL2, tpxh$RWL2$RBL2, tphx$RWL2$RBL2, tplx$RWL2$RBL2, tpxl$RWL2$RBL2);
    if (WWL2==1'b0 && RWL1==1'b0 && RWL2==1'b1 )
       (posedge WWL1 *> (RBL2 -: WBL1)) = (tplh$WWL1$RBL2, tphl$WWL1$RBL2);
    if (WWL2==1'b0 && RWL1==1'b1 && RWL2==1'b0 )
       (posedge WWL1 *> (RBL1 -: WBL1)) = (tplh$WWL1$RBL1, tphl$WWL1$RBL1);
    if (WWL1==1'b0 && RWL1==1'b0 && RWL2==1'b1 )
       (posedge WWL2 *> (RBL2 -: WBL2)) = (tplh$WWL2$RBL2, tphl$WWL2$RBL2);
    if (WWL1==1'b0 && RWL1==1'b1 && RWL2==1'b0 )
       (posedge WWL2 *> (RBL1 -: WBL2)) = (tplh$WWL1$RBL2, tphl$WWL1$RBL2);
    if (WWL1==1'b1 && WWL2==1'b0 && RWL1==1'b1 && RWL2==1'b0 )
       (WBL1 *> RBL1) = (tplh$WBL1$RBL1, tphl$WBL1$RBL1);
    if (WWL1==1'b1 && WWL2==1'b0 && RWL1==1'b0 && RWL2==1'b1 )
       (WBL1 *> RBL2) = (tplh$WBL1$RBL2, tphl$WBL1$RBL2);
    if (WWL1==1'b0 && WWL2==1'b1 && RWL1==1'b1 && RWL2==1'b0 )
       (WBL2 *> RBL1) = (tplh$WBL2$RBL1, tphl$WBL2$RBL1);
    if (WWL1==1'b0 && WWL2==1'b1 && RWL1==1'b0 && RWL2==1'b1 )
       (WBL2 *> RBL2) = (tplh$WBL2$RBL2, tphl$WBL2$RBL2);
    if (WWL2==1'b0 && RWL1==1'b1 && RWL2==1'b1 )
       (posedge WWL1 *> (RBL2 -: WBL1)) = (tplh$WWL1$RBL2, tphl$WWL1$RBL2);
    if (WWL2==1'b0 && RWL1==1'b1 && RWL2==1'b1 )
       (posedge WWL1 *> (RBL1 -: WBL1)) = (tplh$WWL1$RBL1, tphl$WWL1$RBL1);
    if (WWL1==1'b0 && RWL1==1'b1 && RWL2==1'b1 )
       (posedge WWL2 *> (RBL2 -: WBL2)) = (tplh$WWL2$RBL2, tphl$WWL2$RBL2);
    if (WWL1==1'b0 && RWL1==1'b1 && RWL2==1'b1 )
       (posedge WWL2 *> (RBL1 -: WBL2)) = (tplh$WWL1$RBL2, tphl$WWL1$RBL2);
    if (WWL1==1'b1 && WWL2==1'b0 && RWL1==1'b1 && RWL2==1'b1 )
       (WBL1 *> RBL1) = (tplh$WBL1$RBL1, tphl$WBL1$RBL1);
    if (WWL1==1'b1 && WWL2==1'b0 && RWL1==1'b1 && RWL2==1'b1 )
       (WBL1 *> RBL2) = (tplh$WBL1$RBL2, tphl$WBL1$RBL2);
    if (WWL1==1'b0 && WWL2==1'b1 && RWL1==1'b1 && RWL2==1'b1 )
       (WBL2 *> RBL1) = (tplh$WBL2$RBL1, tphl$WBL2$RBL1);
    if (WWL1==1'b0 && WWL2==1'b1 && RWL1==1'b1 && RWL2==1'b1 )
       (WBL2 *> RBL2) = (tplh$WBL2$RBL2, tphl$WBL2$RBL2);
 

  endspecify

endmodule // RF2R2WSX2MA10TR
`endcelldefine
//$Id: rf.genpp,v 1.11 2006/05/18 09:44:11 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module RF2R2WSX1P4MA10TR (RBL1, RBL2, WBL1, WWL1, WBL2, WWL2, RWL1, RWL2);
output RBL1, RBL2;
input WBL1, WWL1, WBL2, WWL2, RWL1, RWL2;
reg NOTIFIER;

   or  I0 (ck, WWL1, WWL2);
   not I1 (ckn, ck);
   udp_wao I2 (wr, WBL1, WBL2, WWL1, WWL2);
   udp_tlatrf I3 (n0, wr, ck, ckn, NOTIFIER);
   not I4 (n1, n0);
   notif1 I5 (RBL1, n1, RWL1);
   notif1 I6 (RBL2, n1, RWL2);

  specify
    // delay parameters
    specparam
      tplh$WBL1$RBL1 = 1.0,
      tphl$WBL1$RBL1 = 1.0,
      tpxh$WBL1$RBL1 = 1.0,
      tphx$WBL1$RBL1 = 1.0,
      tplx$WBL1$RBL1 = 1.0,
      tpxl$WBL1$RBL1 = 1.0,
      tplh$WWL1$RBL1 = 1.0,
      tphl$WWL1$RBL1 = 1.0,
      tpxh$WWL1$RBL1 = 1.0,
      tphx$WWL1$RBL1 = 1.0,
      tplx$WWL1$RBL1 = 1.0,
      tpxl$WWL1$RBL1 = 1.0,
      tplh$WBL2$RBL1 = 1.0,
      tphl$WBL2$RBL1 = 1.0,
      tpxh$WBL2$RBL1 = 1.0,
      tphx$WBL2$RBL1 = 1.0,
      tplx$WBL2$RBL1 = 1.0,
      tpxl$WBL2$RBL1 = 1.0,
      tplh$WWL2$RBL1 = 1.0,
      tphl$WWL2$RBL1 = 1.0,
      tpxh$WWL2$RBL1 = 1.0,
      tphx$WWL2$RBL1 = 1.0,
      tplx$WWL2$RBL1 = 1.0,
      tpxl$WWL2$RBL1 = 1.0,
      tplh$RWL1$RBL1 = 1.0,
      tphl$RWL1$RBL1 = 1.0,
      tpxh$RWL1$RBL1 = 1.0,
      tphx$RWL1$RBL1 = 1.0,
      tplx$RWL1$RBL1 = 1.0,
      tpxl$RWL1$RBL1 = 1.0,
      tplh$RWL2$RBL1 = 1.0,
      tphl$RWL2$RBL1 = 1.0,
      tpxh$RWL2$RBL1 = 1.0,
      tphx$RWL2$RBL1 = 1.0,
      tplx$RWL2$RBL1 = 1.0,
      tpxl$RWL2$RBL1 = 1.0,
      tplh$WBL1$RBL2 = 1.0,
      tphl$WBL1$RBL2 = 1.0,
      tpxh$WBL1$RBL2 = 1.0,
      tphx$WBL1$RBL2 = 1.0,
      tplx$WBL1$RBL2 = 1.0,
      tpxl$WBL1$RBL2 = 1.0,
      tplh$WWL1$RBL2 = 1.0,
      tphl$WWL1$RBL2 = 1.0,
      tpxh$WWL1$RBL2 = 1.0,
      tphx$WWL1$RBL2 = 1.0,
      tplx$WWL1$RBL2 = 1.0,
      tpxl$WWL1$RBL2 = 1.0,
      tplh$WBL2$RBL2 = 1.0,
      tphl$WBL2$RBL2 = 1.0,
      tpxh$WBL2$RBL2 = 1.0,
      tphx$WBL2$RBL2 = 1.0,
      tplx$WBL2$RBL2 = 1.0,
      tpxl$WBL2$RBL2 = 1.0,
      tplh$WWL2$RBL2 = 1.0,
      tphl$WWL2$RBL2 = 1.0,
      tpxh$WWL2$RBL2 = 1.0,
      tphx$WWL2$RBL2 = 1.0,
      tplx$WWL2$RBL2 = 1.0,
      tpxl$WWL2$RBL2 = 1.0,
      tplh$RWL1$RBL2 = 1.0,
      tphl$RWL1$RBL2 = 1.0,
      tpxh$RWL1$RBL2 = 1.0,
      tphx$RWL1$RBL2 = 1.0,
      tplx$RWL1$RBL2 = 1.0,
      tpxl$RWL1$RBL2 = 1.0,
      tplh$RWL2$RBL2 = 1.0,
      tphl$RWL2$RBL2 = 1.0,
      tpxh$RWL2$RBL2 = 1.0,
      tphx$RWL2$RBL2 = 1.0,
      tplx$RWL2$RBL2 = 1.0,
      tpxl$RWL2$RBL2 = 1.0,
    tminpwh$WWL1    = 1.0,
    tperiod$WWL1    = 1.0,
    tminpwh$WWL2    = 1.0,
    tperiod$WWL2    = 1.0,
    tsetup$WWL1$WBL1 = 1.0,
    thold$WWL1$WBL1  = 0.5,
    tsetup$WWL2$WBL2 = 1.0,
    thold$WWL2$WBL2  = 0.5;

      // path delays
 
      // timing checks
      $setuphold(negedge WWL1, posedge WBL1, tsetup$WWL1$WBL1, thold$WWL1$WBL1, NOTIFIER);
      $setuphold(negedge WWL1, negedge WBL1, tsetup$WWL1$WBL1, thold$WWL1$WBL1, NOTIFIER);
      $setuphold(negedge WWL2, posedge WBL2, tsetup$WWL2$WBL2, thold$WWL2$WBL2, NOTIFIER);
      $setuphold(negedge WWL2, negedge WBL2, tsetup$WWL2$WBL2, thold$WWL2$WBL2, NOTIFIER);
      $width(posedge WWL1, tminpwh$WWL1, 0, NOTIFIER);
      $period(posedge WWL1, tperiod$WWL1, NOTIFIER);
      $width(posedge WWL2, tminpwh$WWL2, 0, NOTIFIER);
      $period(posedge WWL2, tperiod$WWL2, NOTIFIER);
    if (WWL1==1'b0 && WWL2==1'b0 && RWL2==1'b0 )
       (RWL1 *> RBL1) = (tplh$RWL1$RBL1, tphl$RWL1$RBL1, tpxh$RWL1$RBL1, tphx$RWL1$RBL1, tplx$RWL1$RBL1, tpxl$RWL1$RBL1);
    if (WWL1==1'b0 && WWL2==1'b0 && RWL1==1'b0 )
       (RWL2 *> RBL2) = (tplh$RWL2$RBL2, tphl$RWL2$RBL2, tpxh$RWL2$RBL2, tphx$RWL2$RBL2, tplx$RWL2$RBL2, tpxl$RWL2$RBL2);
    if (WWL1==1'b0 && WWL2==1'b0 && RWL2==1'b1 )
       (RWL1 *> RBL1) = (tplh$RWL1$RBL1, tphl$RWL1$RBL1, tpxh$RWL1$RBL1, tphx$RWL1$RBL1, tplx$RWL1$RBL1, tpxl$RWL1$RBL1);
    if (WWL1==1'b0 && WWL2==1'b0 && RWL1==1'b1 )
       (RWL2 *> RBL2) = (tplh$RWL2$RBL2, tphl$RWL2$RBL2, tpxh$RWL2$RBL2, tphx$RWL2$RBL2, tplx$RWL2$RBL2, tpxl$RWL2$RBL2);
    if (WWL1==1'b0 && WWL2==1'b1 && RWL2==1'b0 )
       (RWL1 *> RBL1) = (tplh$RWL1$RBL1, tphl$RWL1$RBL1, tpxh$RWL1$RBL1, tphx$RWL1$RBL1, tplx$RWL1$RBL1, tpxl$RWL1$RBL1);
    if (WWL1==1'b0 && WWL2==1'b1 && RWL1==1'b0 )
       (RWL2 *> RBL2) = (tplh$RWL2$RBL2, tphl$RWL2$RBL2, tpxh$RWL2$RBL2, tphx$RWL2$RBL2, tplx$RWL2$RBL2, tpxl$RWL2$RBL2);
    if (WWL1==1'b0 && WWL2==1'b1 && RWL2==1'b1 )
       (RWL1 *> RBL1) = (tplh$RWL1$RBL1, tphl$RWL1$RBL1, tpxh$RWL1$RBL1, tphx$RWL1$RBL1, tplx$RWL1$RBL1, tpxl$RWL1$RBL1);
    if (WWL1==1'b0 && WWL2==1'b1 && RWL1==1'b1 )
       (RWL2 *> RBL2) = (tplh$RWL2$RBL2, tphl$RWL2$RBL2, tpxh$RWL2$RBL2, tphx$RWL2$RBL2, tplx$RWL2$RBL2, tpxl$RWL2$RBL2);
    if (WWL1==1'b1 && WWL2==1'b0 && RWL2==1'b0 )
       (RWL1 *> RBL1) = (tplh$RWL1$RBL1, tphl$RWL1$RBL1, tpxh$RWL1$RBL1, tphx$RWL1$RBL1, tplx$RWL1$RBL1, tpxl$RWL1$RBL1);
    if (WWL1==1'b1 && WWL2==1'b0 && RWL1==1'b0 )
       (RWL2 *> RBL2) = (tplh$RWL2$RBL2, tphl$RWL2$RBL2, tpxh$RWL2$RBL2, tphx$RWL2$RBL2, tplx$RWL2$RBL2, tpxl$RWL2$RBL2);
    if (WWL1==1'b1 && WWL2==1'b0 && RWL2==1'b1 )
       (RWL1 *> RBL1) = (tplh$RWL1$RBL1, tphl$RWL1$RBL1, tpxh$RWL1$RBL1, tphx$RWL1$RBL1, tplx$RWL1$RBL1, tpxl$RWL1$RBL1);
    if (WWL1==1'b1 && WWL2==1'b0 && RWL1==1'b1 )
       (RWL2 *> RBL2) = (tplh$RWL2$RBL2, tphl$RWL2$RBL2, tpxh$RWL2$RBL2, tphx$RWL2$RBL2, tplx$RWL2$RBL2, tpxl$RWL2$RBL2);
    if (WWL1==1'b1 && WWL2==1'b1 && RWL2==1'b0 )
       (RWL1 *> RBL1) = (tplh$RWL1$RBL1, tphl$RWL1$RBL1, tpxh$RWL1$RBL1, tphx$RWL1$RBL1, tplx$RWL1$RBL1, tpxl$RWL1$RBL1);
    if (WWL1==1'b1 && WWL2==1'b1 && RWL1==1'b0 )
       (RWL2 *> RBL2) = (tplh$RWL2$RBL2, tphl$RWL2$RBL2, tpxh$RWL2$RBL2, tphx$RWL2$RBL2, tplx$RWL2$RBL2, tpxl$RWL2$RBL2);
    if (WWL1==1'b1 && WWL2==1'b1 && RWL2==1'b1 )
       (RWL1 *> RBL1) = (tplh$RWL1$RBL1, tphl$RWL1$RBL1, tpxh$RWL1$RBL1, tphx$RWL1$RBL1, tplx$RWL1$RBL1, tpxl$RWL1$RBL1);
    if (WWL1==1'b1 && WWL2==1'b1 && RWL1==1'b1 )
       (RWL2 *> RBL2) = (tplh$RWL2$RBL2, tphl$RWL2$RBL2, tpxh$RWL2$RBL2, tphx$RWL2$RBL2, tplx$RWL2$RBL2, tpxl$RWL2$RBL2);
    if (WWL2==1'b0 && RWL1==1'b0 && RWL2==1'b1 )
       (posedge WWL1 *> (RBL2 -: WBL1)) = (tplh$WWL1$RBL2, tphl$WWL1$RBL2);
    if (WWL2==1'b0 && RWL1==1'b1 && RWL2==1'b0 )
       (posedge WWL1 *> (RBL1 -: WBL1)) = (tplh$WWL1$RBL1, tphl$WWL1$RBL1);
    if (WWL1==1'b0 && RWL1==1'b0 && RWL2==1'b1 )
       (posedge WWL2 *> (RBL2 -: WBL2)) = (tplh$WWL2$RBL2, tphl$WWL2$RBL2);
    if (WWL1==1'b0 && RWL1==1'b1 && RWL2==1'b0 )
       (posedge WWL2 *> (RBL1 -: WBL2)) = (tplh$WWL1$RBL2, tphl$WWL1$RBL2);
    if (WWL1==1'b1 && WWL2==1'b0 && RWL1==1'b1 && RWL2==1'b0 )
       (WBL1 *> RBL1) = (tplh$WBL1$RBL1, tphl$WBL1$RBL1);
    if (WWL1==1'b1 && WWL2==1'b0 && RWL1==1'b0 && RWL2==1'b1 )
       (WBL1 *> RBL2) = (tplh$WBL1$RBL2, tphl$WBL1$RBL2);
    if (WWL1==1'b0 && WWL2==1'b1 && RWL1==1'b1 && RWL2==1'b0 )
       (WBL2 *> RBL1) = (tplh$WBL2$RBL1, tphl$WBL2$RBL1);
    if (WWL1==1'b0 && WWL2==1'b1 && RWL1==1'b0 && RWL2==1'b1 )
       (WBL2 *> RBL2) = (tplh$WBL2$RBL2, tphl$WBL2$RBL2);
    if (WWL2==1'b0 && RWL1==1'b1 && RWL2==1'b1 )
       (posedge WWL1 *> (RBL2 -: WBL1)) = (tplh$WWL1$RBL2, tphl$WWL1$RBL2);
    if (WWL2==1'b0 && RWL1==1'b1 && RWL2==1'b1 )
       (posedge WWL1 *> (RBL1 -: WBL1)) = (tplh$WWL1$RBL1, tphl$WWL1$RBL1);
    if (WWL1==1'b0 && RWL1==1'b1 && RWL2==1'b1 )
       (posedge WWL2 *> (RBL2 -: WBL2)) = (tplh$WWL2$RBL2, tphl$WWL2$RBL2);
    if (WWL1==1'b0 && RWL1==1'b1 && RWL2==1'b1 )
       (posedge WWL2 *> (RBL1 -: WBL2)) = (tplh$WWL1$RBL2, tphl$WWL1$RBL2);
    if (WWL1==1'b1 && WWL2==1'b0 && RWL1==1'b1 && RWL2==1'b1 )
       (WBL1 *> RBL1) = (tplh$WBL1$RBL1, tphl$WBL1$RBL1);
    if (WWL1==1'b1 && WWL2==1'b0 && RWL1==1'b1 && RWL2==1'b1 )
       (WBL1 *> RBL2) = (tplh$WBL1$RBL2, tphl$WBL1$RBL2);
    if (WWL1==1'b0 && WWL2==1'b1 && RWL1==1'b1 && RWL2==1'b1 )
       (WBL2 *> RBL1) = (tplh$WBL2$RBL1, tphl$WBL2$RBL1);
    if (WWL1==1'b0 && WWL2==1'b1 && RWL1==1'b1 && RWL2==1'b1 )
       (WBL2 *> RBL2) = (tplh$WBL2$RBL2, tphl$WBL2$RBL2);
 

  endspecify

endmodule // RF2R2WSX1P4MA10TR
`endcelldefine
//$Id: rf.genpp,v 1.11 2006/05/18 09:44:11 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module RF2R2WSX1MA10TR (RBL1, RBL2, WBL1, WWL1, WBL2, WWL2, RWL1, RWL2);
output RBL1, RBL2;
input WBL1, WWL1, WBL2, WWL2, RWL1, RWL2;
reg NOTIFIER;

   or  I0 (ck, WWL1, WWL2);
   not I1 (ckn, ck);
   udp_wao I2 (wr, WBL1, WBL2, WWL1, WWL2);
   udp_tlatrf I3 (n0, wr, ck, ckn, NOTIFIER);
   not I4 (n1, n0);
   notif1 I5 (RBL1, n1, RWL1);
   notif1 I6 (RBL2, n1, RWL2);

  specify
    // delay parameters
    specparam
      tplh$WBL1$RBL1 = 1.0,
      tphl$WBL1$RBL1 = 1.0,
      tpxh$WBL1$RBL1 = 1.0,
      tphx$WBL1$RBL1 = 1.0,
      tplx$WBL1$RBL1 = 1.0,
      tpxl$WBL1$RBL1 = 1.0,
      tplh$WWL1$RBL1 = 1.0,
      tphl$WWL1$RBL1 = 1.0,
      tpxh$WWL1$RBL1 = 1.0,
      tphx$WWL1$RBL1 = 1.0,
      tplx$WWL1$RBL1 = 1.0,
      tpxl$WWL1$RBL1 = 1.0,
      tplh$WBL2$RBL1 = 1.0,
      tphl$WBL2$RBL1 = 1.0,
      tpxh$WBL2$RBL1 = 1.0,
      tphx$WBL2$RBL1 = 1.0,
      tplx$WBL2$RBL1 = 1.0,
      tpxl$WBL2$RBL1 = 1.0,
      tplh$WWL2$RBL1 = 1.0,
      tphl$WWL2$RBL1 = 1.0,
      tpxh$WWL2$RBL1 = 1.0,
      tphx$WWL2$RBL1 = 1.0,
      tplx$WWL2$RBL1 = 1.0,
      tpxl$WWL2$RBL1 = 1.0,
      tplh$RWL1$RBL1 = 1.0,
      tphl$RWL1$RBL1 = 1.0,
      tpxh$RWL1$RBL1 = 1.0,
      tphx$RWL1$RBL1 = 1.0,
      tplx$RWL1$RBL1 = 1.0,
      tpxl$RWL1$RBL1 = 1.0,
      tplh$RWL2$RBL1 = 1.0,
      tphl$RWL2$RBL1 = 1.0,
      tpxh$RWL2$RBL1 = 1.0,
      tphx$RWL2$RBL1 = 1.0,
      tplx$RWL2$RBL1 = 1.0,
      tpxl$RWL2$RBL1 = 1.0,
      tplh$WBL1$RBL2 = 1.0,
      tphl$WBL1$RBL2 = 1.0,
      tpxh$WBL1$RBL2 = 1.0,
      tphx$WBL1$RBL2 = 1.0,
      tplx$WBL1$RBL2 = 1.0,
      tpxl$WBL1$RBL2 = 1.0,
      tplh$WWL1$RBL2 = 1.0,
      tphl$WWL1$RBL2 = 1.0,
      tpxh$WWL1$RBL2 = 1.0,
      tphx$WWL1$RBL2 = 1.0,
      tplx$WWL1$RBL2 = 1.0,
      tpxl$WWL1$RBL2 = 1.0,
      tplh$WBL2$RBL2 = 1.0,
      tphl$WBL2$RBL2 = 1.0,
      tpxh$WBL2$RBL2 = 1.0,
      tphx$WBL2$RBL2 = 1.0,
      tplx$WBL2$RBL2 = 1.0,
      tpxl$WBL2$RBL2 = 1.0,
      tplh$WWL2$RBL2 = 1.0,
      tphl$WWL2$RBL2 = 1.0,
      tpxh$WWL2$RBL2 = 1.0,
      tphx$WWL2$RBL2 = 1.0,
      tplx$WWL2$RBL2 = 1.0,
      tpxl$WWL2$RBL2 = 1.0,
      tplh$RWL1$RBL2 = 1.0,
      tphl$RWL1$RBL2 = 1.0,
      tpxh$RWL1$RBL2 = 1.0,
      tphx$RWL1$RBL2 = 1.0,
      tplx$RWL1$RBL2 = 1.0,
      tpxl$RWL1$RBL2 = 1.0,
      tplh$RWL2$RBL2 = 1.0,
      tphl$RWL2$RBL2 = 1.0,
      tpxh$RWL2$RBL2 = 1.0,
      tphx$RWL2$RBL2 = 1.0,
      tplx$RWL2$RBL2 = 1.0,
      tpxl$RWL2$RBL2 = 1.0,
    tminpwh$WWL1    = 1.0,
    tperiod$WWL1    = 1.0,
    tminpwh$WWL2    = 1.0,
    tperiod$WWL2    = 1.0,
    tsetup$WWL1$WBL1 = 1.0,
    thold$WWL1$WBL1  = 0.5,
    tsetup$WWL2$WBL2 = 1.0,
    thold$WWL2$WBL2  = 0.5;

      // path delays
 
      // timing checks
      $setuphold(negedge WWL1, posedge WBL1, tsetup$WWL1$WBL1, thold$WWL1$WBL1, NOTIFIER);
      $setuphold(negedge WWL1, negedge WBL1, tsetup$WWL1$WBL1, thold$WWL1$WBL1, NOTIFIER);
      $setuphold(negedge WWL2, posedge WBL2, tsetup$WWL2$WBL2, thold$WWL2$WBL2, NOTIFIER);
      $setuphold(negedge WWL2, negedge WBL2, tsetup$WWL2$WBL2, thold$WWL2$WBL2, NOTIFIER);
      $width(posedge WWL1, tminpwh$WWL1, 0, NOTIFIER);
      $period(posedge WWL1, tperiod$WWL1, NOTIFIER);
      $width(posedge WWL2, tminpwh$WWL2, 0, NOTIFIER);
      $period(posedge WWL2, tperiod$WWL2, NOTIFIER);
    if (WWL1==1'b0 && WWL2==1'b0 && RWL2==1'b0 )
       (RWL1 *> RBL1) = (tplh$RWL1$RBL1, tphl$RWL1$RBL1, tpxh$RWL1$RBL1, tphx$RWL1$RBL1, tplx$RWL1$RBL1, tpxl$RWL1$RBL1);
    if (WWL1==1'b0 && WWL2==1'b0 && RWL1==1'b0 )
       (RWL2 *> RBL2) = (tplh$RWL2$RBL2, tphl$RWL2$RBL2, tpxh$RWL2$RBL2, tphx$RWL2$RBL2, tplx$RWL2$RBL2, tpxl$RWL2$RBL2);
    if (WWL1==1'b0 && WWL2==1'b0 && RWL2==1'b1 )
       (RWL1 *> RBL1) = (tplh$RWL1$RBL1, tphl$RWL1$RBL1, tpxh$RWL1$RBL1, tphx$RWL1$RBL1, tplx$RWL1$RBL1, tpxl$RWL1$RBL1);
    if (WWL1==1'b0 && WWL2==1'b0 && RWL1==1'b1 )
       (RWL2 *> RBL2) = (tplh$RWL2$RBL2, tphl$RWL2$RBL2, tpxh$RWL2$RBL2, tphx$RWL2$RBL2, tplx$RWL2$RBL2, tpxl$RWL2$RBL2);
    if (WWL1==1'b0 && WWL2==1'b1 && RWL2==1'b0 )
       (RWL1 *> RBL1) = (tplh$RWL1$RBL1, tphl$RWL1$RBL1, tpxh$RWL1$RBL1, tphx$RWL1$RBL1, tplx$RWL1$RBL1, tpxl$RWL1$RBL1);
    if (WWL1==1'b0 && WWL2==1'b1 && RWL1==1'b0 )
       (RWL2 *> RBL2) = (tplh$RWL2$RBL2, tphl$RWL2$RBL2, tpxh$RWL2$RBL2, tphx$RWL2$RBL2, tplx$RWL2$RBL2, tpxl$RWL2$RBL2);
    if (WWL1==1'b0 && WWL2==1'b1 && RWL2==1'b1 )
       (RWL1 *> RBL1) = (tplh$RWL1$RBL1, tphl$RWL1$RBL1, tpxh$RWL1$RBL1, tphx$RWL1$RBL1, tplx$RWL1$RBL1, tpxl$RWL1$RBL1);
    if (WWL1==1'b0 && WWL2==1'b1 && RWL1==1'b1 )
       (RWL2 *> RBL2) = (tplh$RWL2$RBL2, tphl$RWL2$RBL2, tpxh$RWL2$RBL2, tphx$RWL2$RBL2, tplx$RWL2$RBL2, tpxl$RWL2$RBL2);
    if (WWL1==1'b1 && WWL2==1'b0 && RWL2==1'b0 )
       (RWL1 *> RBL1) = (tplh$RWL1$RBL1, tphl$RWL1$RBL1, tpxh$RWL1$RBL1, tphx$RWL1$RBL1, tplx$RWL1$RBL1, tpxl$RWL1$RBL1);
    if (WWL1==1'b1 && WWL2==1'b0 && RWL1==1'b0 )
       (RWL2 *> RBL2) = (tplh$RWL2$RBL2, tphl$RWL2$RBL2, tpxh$RWL2$RBL2, tphx$RWL2$RBL2, tplx$RWL2$RBL2, tpxl$RWL2$RBL2);
    if (WWL1==1'b1 && WWL2==1'b0 && RWL2==1'b1 )
       (RWL1 *> RBL1) = (tplh$RWL1$RBL1, tphl$RWL1$RBL1, tpxh$RWL1$RBL1, tphx$RWL1$RBL1, tplx$RWL1$RBL1, tpxl$RWL1$RBL1);
    if (WWL1==1'b1 && WWL2==1'b0 && RWL1==1'b1 )
       (RWL2 *> RBL2) = (tplh$RWL2$RBL2, tphl$RWL2$RBL2, tpxh$RWL2$RBL2, tphx$RWL2$RBL2, tplx$RWL2$RBL2, tpxl$RWL2$RBL2);
    if (WWL1==1'b1 && WWL2==1'b1 && RWL2==1'b0 )
       (RWL1 *> RBL1) = (tplh$RWL1$RBL1, tphl$RWL1$RBL1, tpxh$RWL1$RBL1, tphx$RWL1$RBL1, tplx$RWL1$RBL1, tpxl$RWL1$RBL1);
    if (WWL1==1'b1 && WWL2==1'b1 && RWL1==1'b0 )
       (RWL2 *> RBL2) = (tplh$RWL2$RBL2, tphl$RWL2$RBL2, tpxh$RWL2$RBL2, tphx$RWL2$RBL2, tplx$RWL2$RBL2, tpxl$RWL2$RBL2);
    if (WWL1==1'b1 && WWL2==1'b1 && RWL2==1'b1 )
       (RWL1 *> RBL1) = (tplh$RWL1$RBL1, tphl$RWL1$RBL1, tpxh$RWL1$RBL1, tphx$RWL1$RBL1, tplx$RWL1$RBL1, tpxl$RWL1$RBL1);
    if (WWL1==1'b1 && WWL2==1'b1 && RWL1==1'b1 )
       (RWL2 *> RBL2) = (tplh$RWL2$RBL2, tphl$RWL2$RBL2, tpxh$RWL2$RBL2, tphx$RWL2$RBL2, tplx$RWL2$RBL2, tpxl$RWL2$RBL2);
    if (WWL2==1'b0 && RWL1==1'b0 && RWL2==1'b1 )
       (posedge WWL1 *> (RBL2 -: WBL1)) = (tplh$WWL1$RBL2, tphl$WWL1$RBL2);
    if (WWL2==1'b0 && RWL1==1'b1 && RWL2==1'b0 )
       (posedge WWL1 *> (RBL1 -: WBL1)) = (tplh$WWL1$RBL1, tphl$WWL1$RBL1);
    if (WWL1==1'b0 && RWL1==1'b0 && RWL2==1'b1 )
       (posedge WWL2 *> (RBL2 -: WBL2)) = (tplh$WWL2$RBL2, tphl$WWL2$RBL2);
    if (WWL1==1'b0 && RWL1==1'b1 && RWL2==1'b0 )
       (posedge WWL2 *> (RBL1 -: WBL2)) = (tplh$WWL1$RBL2, tphl$WWL1$RBL2);
    if (WWL1==1'b1 && WWL2==1'b0 && RWL1==1'b1 && RWL2==1'b0 )
       (WBL1 *> RBL1) = (tplh$WBL1$RBL1, tphl$WBL1$RBL1);
    if (WWL1==1'b1 && WWL2==1'b0 && RWL1==1'b0 && RWL2==1'b1 )
       (WBL1 *> RBL2) = (tplh$WBL1$RBL2, tphl$WBL1$RBL2);
    if (WWL1==1'b0 && WWL2==1'b1 && RWL1==1'b1 && RWL2==1'b0 )
       (WBL2 *> RBL1) = (tplh$WBL2$RBL1, tphl$WBL2$RBL1);
    if (WWL1==1'b0 && WWL2==1'b1 && RWL1==1'b0 && RWL2==1'b1 )
       (WBL2 *> RBL2) = (tplh$WBL2$RBL2, tphl$WBL2$RBL2);
    if (WWL2==1'b0 && RWL1==1'b1 && RWL2==1'b1 )
       (posedge WWL1 *> (RBL2 -: WBL1)) = (tplh$WWL1$RBL2, tphl$WWL1$RBL2);
    if (WWL2==1'b0 && RWL1==1'b1 && RWL2==1'b1 )
       (posedge WWL1 *> (RBL1 -: WBL1)) = (tplh$WWL1$RBL1, tphl$WWL1$RBL1);
    if (WWL1==1'b0 && RWL1==1'b1 && RWL2==1'b1 )
       (posedge WWL2 *> (RBL2 -: WBL2)) = (tplh$WWL2$RBL2, tphl$WWL2$RBL2);
    if (WWL1==1'b0 && RWL1==1'b1 && RWL2==1'b1 )
       (posedge WWL2 *> (RBL1 -: WBL2)) = (tplh$WWL1$RBL2, tphl$WWL1$RBL2);
    if (WWL1==1'b1 && WWL2==1'b0 && RWL1==1'b1 && RWL2==1'b1 )
       (WBL1 *> RBL1) = (tplh$WBL1$RBL1, tphl$WBL1$RBL1);
    if (WWL1==1'b1 && WWL2==1'b0 && RWL1==1'b1 && RWL2==1'b1 )
       (WBL1 *> RBL2) = (tplh$WBL1$RBL2, tphl$WBL1$RBL2);
    if (WWL1==1'b0 && WWL2==1'b1 && RWL1==1'b1 && RWL2==1'b1 )
       (WBL2 *> RBL1) = (tplh$WBL2$RBL1, tphl$WBL2$RBL1);
    if (WWL1==1'b0 && WWL2==1'b1 && RWL1==1'b1 && RWL2==1'b1 )
       (WBL2 *> RBL2) = (tplh$WBL2$RBL2, tphl$WBL2$RBL2);
 

  endspecify

endmodule // RF2R2WSX1MA10TR
`endcelldefine
//$Id: rf.genpp,v 1.11 2006/05/18 09:44:11 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module RF2R1WSX2MA10TR (RBL1, RBL2, WBL, WWL, RWL1, RWL2);
output RBL1, RBL2;
input WBL, WWL, RWL1, RWL2;
reg NOTIFIER;

   not        I0 (WWLN, WWL);
   not        I1 (R1WN, RWL1);
   not        I2 (RWL2N, RWL2);
   udp_tlatrf I3 (n0, WBL, WWL, WWLN, NOTIFIER);
   bufif1     I4 (RBL1, n0, n2);
   bufif1     I5 (RBL2, n0, n3);
   udp_outrf  I6 (n2, n0, R1WN, RWL1);
   udp_outrf  I7 (n3, n0, RWL2N, RWL2);

  specify
    // delay parameters
    specparam
      tplh$WBL$RBL1 = 1.0,
      tphl$WBL$RBL1 = 1.0,
      tpxh$WBL$RBL1 = 1.0,
      tphx$WBL$RBL1 = 1.0,
      tplx$WBL$RBL1 = 1.0,
      tpxl$WBL$RBL1 = 1.0,
      tplh$WWL$RBL1 = 1.0,
      tphl$WWL$RBL1 = 1.0,
      tpxh$WWL$RBL1 = 1.0,
      tphx$WWL$RBL1 = 1.0,
      tplx$WWL$RBL1 = 1.0,
      tpxl$WWL$RBL1 = 1.0,
      tplh$RWL1$RBL1 = 1.0,
      tphl$RWL1$RBL1 = 1.0,
      tpxh$RWL1$RBL1 = 1.0,
      tphx$RWL1$RBL1 = 1.0,
      tplx$RWL1$RBL1 = 1.0,
      tpxl$RWL1$RBL1 = 1.0,
      tplh$RWL2$RBL1 = 1.0,
      tphl$RWL2$RBL1 = 1.0,
      tpxh$RWL2$RBL1 = 1.0,
      tphx$RWL2$RBL1 = 1.0,
      tplx$RWL2$RBL1 = 1.0,
      tpxl$RWL2$RBL1 = 1.0,
      tplh$WBL$RBL2 = 1.0,
      tphl$WBL$RBL2 = 1.0,
      tpxh$WBL$RBL2 = 1.0,
      tphx$WBL$RBL2 = 1.0,
      tplx$WBL$RBL2 = 1.0,
      tpxl$WBL$RBL2 = 1.0,
      tplh$WWL$RBL2 = 1.0,
      tphl$WWL$RBL2 = 1.0,
      tpxh$WWL$RBL2 = 1.0,
      tphx$WWL$RBL2 = 1.0,
      tplx$WWL$RBL2 = 1.0,
      tpxl$WWL$RBL2 = 1.0,
      tplh$RWL1$RBL2 = 1.0,
      tphl$RWL1$RBL2 = 1.0,
      tpxh$RWL1$RBL2 = 1.0,
      tphx$RWL1$RBL2 = 1.0,
      tplx$RWL1$RBL2 = 1.0,
      tpxl$RWL1$RBL2 = 1.0,
      tplh$RWL2$RBL2 = 1.0,
      tphl$RWL2$RBL2 = 1.0,
      tpxh$RWL2$RBL2 = 1.0,
      tphx$RWL2$RBL2 = 1.0,
      tplx$RWL2$RBL2 = 1.0,
      tpxl$RWL2$RBL2 = 1.0,
    tminpwh$WWL    = 1.0,
    tperiod$WWL    = 1.0,
    tsetup$WWL$WBL = 1.0,
    thold$WWL$WBL  = 0.5;

      // path delays
      ( WWL *> RBL1) = (tplh$WWL$RBL1, tphl$WWL$RBL1);
      ( WWL *> RBL2) = (tplh$WWL$RBL2, tphl$WWL$RBL2);
 
      // timing checks
      $width(posedge WWL, tminpwh$WWL, 0, NOTIFIER);
      $period(posedge WWL, tperiod$WWL, NOTIFIER);
      $setuphold(negedge WWL, posedge WBL, tsetup$WWL$WBL, thold$WWL$WBL, NOTIFIER);
      $setuphold(negedge WWL, negedge WBL, tsetup$WWL$WBL, thold$WWL$WBL, NOTIFIER);
    if (WBL==1'b0 && WWL==1'b0 && RWL2==1'b0 )
       (RWL1 *> RBL1) = (tplh$RWL1$RBL1, tphl$RWL1$RBL1, tpxh$RWL1$RBL1, tphx$RWL1$RBL1, tplx$RWL1$RBL1, tpxl$RWL1$RBL1);
    if (WBL==1'b0 && WWL==1'b0 && RWL1==1'b0 )
       (RWL2 *> RBL2) = (tplh$RWL2$RBL2, tphl$RWL2$RBL2, tpxh$RWL2$RBL2, tphx$RWL2$RBL2, tplx$RWL2$RBL2, tpxl$RWL2$RBL2);
    if (WBL==1'b0 && WWL==1'b0 && RWL2==1'b1 )
       (RWL1 *> RBL1) = (tplh$RWL1$RBL1, tphl$RWL1$RBL1, tpxh$RWL1$RBL1, tphx$RWL1$RBL1, tplx$RWL1$RBL1, tpxl$RWL1$RBL1);
    if (WBL==1'b0 && WWL==1'b0 && RWL1==1'b1 )
       (RWL2 *> RBL2) = (tplh$RWL2$RBL2, tphl$RWL2$RBL2, tpxh$RWL2$RBL2, tphx$RWL2$RBL2, tplx$RWL2$RBL2, tpxl$RWL2$RBL2);
    if (WBL==1'b1 && WWL==1'b0 && RWL2==1'b0 )
       (RWL1 *> RBL1) = (tplh$RWL1$RBL1, tphl$RWL1$RBL1, tpxh$RWL1$RBL1, tphx$RWL1$RBL1, tplx$RWL1$RBL1, tpxl$RWL1$RBL1);
    if (WBL==1'b1 && WWL==1'b0 && RWL1==1'b0 )
       (RWL2 *> RBL2) = (tplh$RWL2$RBL2, tphl$RWL2$RBL2, tpxh$RWL2$RBL2, tphx$RWL2$RBL2, tplx$RWL2$RBL2, tpxl$RWL2$RBL2);
    if (WBL==1'b1 && WWL==1'b0 && RWL2==1'b1 )
       (RWL1 *> RBL1) = (tplh$RWL1$RBL1, tphl$RWL1$RBL1, tpxh$RWL1$RBL1, tphx$RWL1$RBL1, tplx$RWL1$RBL1, tpxl$RWL1$RBL1);
    if (WBL==1'b1 && WWL==1'b0 && RWL1==1'b1 )
       (RWL2 *> RBL2) = (tplh$RWL2$RBL2, tphl$RWL2$RBL2, tpxh$RWL2$RBL2, tphx$RWL2$RBL2, tplx$RWL2$RBL2, tpxl$RWL2$RBL2);
    if (WWL==1'b1 && RWL2==1'b0 )
       (RWL1 *> RBL1) = (tplh$RWL1$RBL1, tphl$RWL1$RBL1, tpxh$RWL1$RBL1, tphx$RWL1$RBL1, tplx$RWL1$RBL1, tpxl$RWL1$RBL1);
    if (WWL==1'b1 && RWL1==1'b0 )
       (RWL2 *> RBL2) = (tplh$RWL2$RBL2, tphl$RWL2$RBL2, tpxh$RWL2$RBL2, tphx$RWL2$RBL2, tplx$RWL2$RBL2, tpxl$RWL2$RBL2);
    if (WWL==1'b1 &&  RWL2==1'b0 )
       (WBL *> RBL1) = (tplh$WBL$RBL1, tphl$WBL$RBL1);
    if (WWL==1'b1 && RWL1==1'b0 )
       (WBL *> RBL2) = (tplh$WBL$RBL2, tphl$WBL$RBL2);
    if (WWL==1'b1 && RWL2==1'b1 )
       (RWL1 *> RBL1) = (tplh$RWL1$RBL1, tphl$RWL1$RBL1, tpxh$RWL1$RBL1, tphx$RWL1$RBL1, tplx$RWL1$RBL1, tpxl$RWL1$RBL1);
    if (WWL==1'b1 && RWL1==1'b1 )
       (RWL2 *> RBL2) = (tplh$RWL2$RBL2, tphl$RWL2$RBL2, tpxh$RWL2$RBL2, tphx$RWL2$RBL2, tplx$RWL2$RBL2, tpxl$RWL2$RBL2);
    if (WWL==1'b1 &&  RWL2==1'b1 )
       (WBL *> RBL1) = (tplh$WBL$RBL1, tphl$WBL$RBL1);
    if (WWL==1'b1 && RWL1==1'b1 )
       (WBL *> RBL2) = (tplh$WBL$RBL2, tphl$WBL$RBL2);
 

  endspecify

endmodule // RF2R1WSX2MA10TR
`endcelldefine
//$Id: rf.genpp,v 1.11 2006/05/18 09:44:11 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module RF2R1WSX1P4MA10TR (RBL1, RBL2, WBL, WWL, RWL1, RWL2);
output RBL1, RBL2;
input WBL, WWL, RWL1, RWL2;
reg NOTIFIER;

   not        I0 (WWLN, WWL);
   not        I1 (R1WN, RWL1);
   not        I2 (RWL2N, RWL2);
   udp_tlatrf I3 (n0, WBL, WWL, WWLN, NOTIFIER);
   bufif1     I4 (RBL1, n0, n2);
   bufif1     I5 (RBL2, n0, n3);
   udp_outrf  I6 (n2, n0, R1WN, RWL1);
   udp_outrf  I7 (n3, n0, RWL2N, RWL2);

  specify
    // delay parameters
    specparam
      tplh$WBL$RBL1 = 1.0,
      tphl$WBL$RBL1 = 1.0,
      tpxh$WBL$RBL1 = 1.0,
      tphx$WBL$RBL1 = 1.0,
      tplx$WBL$RBL1 = 1.0,
      tpxl$WBL$RBL1 = 1.0,
      tplh$WWL$RBL1 = 1.0,
      tphl$WWL$RBL1 = 1.0,
      tpxh$WWL$RBL1 = 1.0,
      tphx$WWL$RBL1 = 1.0,
      tplx$WWL$RBL1 = 1.0,
      tpxl$WWL$RBL1 = 1.0,
      tplh$RWL1$RBL1 = 1.0,
      tphl$RWL1$RBL1 = 1.0,
      tpxh$RWL1$RBL1 = 1.0,
      tphx$RWL1$RBL1 = 1.0,
      tplx$RWL1$RBL1 = 1.0,
      tpxl$RWL1$RBL1 = 1.0,
      tplh$RWL2$RBL1 = 1.0,
      tphl$RWL2$RBL1 = 1.0,
      tpxh$RWL2$RBL1 = 1.0,
      tphx$RWL2$RBL1 = 1.0,
      tplx$RWL2$RBL1 = 1.0,
      tpxl$RWL2$RBL1 = 1.0,
      tplh$WBL$RBL2 = 1.0,
      tphl$WBL$RBL2 = 1.0,
      tpxh$WBL$RBL2 = 1.0,
      tphx$WBL$RBL2 = 1.0,
      tplx$WBL$RBL2 = 1.0,
      tpxl$WBL$RBL2 = 1.0,
      tplh$WWL$RBL2 = 1.0,
      tphl$WWL$RBL2 = 1.0,
      tpxh$WWL$RBL2 = 1.0,
      tphx$WWL$RBL2 = 1.0,
      tplx$WWL$RBL2 = 1.0,
      tpxl$WWL$RBL2 = 1.0,
      tplh$RWL1$RBL2 = 1.0,
      tphl$RWL1$RBL2 = 1.0,
      tpxh$RWL1$RBL2 = 1.0,
      tphx$RWL1$RBL2 = 1.0,
      tplx$RWL1$RBL2 = 1.0,
      tpxl$RWL1$RBL2 = 1.0,
      tplh$RWL2$RBL2 = 1.0,
      tphl$RWL2$RBL2 = 1.0,
      tpxh$RWL2$RBL2 = 1.0,
      tphx$RWL2$RBL2 = 1.0,
      tplx$RWL2$RBL2 = 1.0,
      tpxl$RWL2$RBL2 = 1.0,
    tminpwh$WWL    = 1.0,
    tperiod$WWL    = 1.0,
    tsetup$WWL$WBL = 1.0,
    thold$WWL$WBL  = 0.5;

      // path delays
      ( WWL *> RBL1) = (tplh$WWL$RBL1, tphl$WWL$RBL1);
      ( WWL *> RBL2) = (tplh$WWL$RBL2, tphl$WWL$RBL2);
 
      // timing checks
      $width(posedge WWL, tminpwh$WWL, 0, NOTIFIER);
      $period(posedge WWL, tperiod$WWL, NOTIFIER);
      $setuphold(negedge WWL, posedge WBL, tsetup$WWL$WBL, thold$WWL$WBL, NOTIFIER);
      $setuphold(negedge WWL, negedge WBL, tsetup$WWL$WBL, thold$WWL$WBL, NOTIFIER);
    if (WBL==1'b0 && WWL==1'b0 && RWL2==1'b0 )
       (RWL1 *> RBL1) = (tplh$RWL1$RBL1, tphl$RWL1$RBL1, tpxh$RWL1$RBL1, tphx$RWL1$RBL1, tplx$RWL1$RBL1, tpxl$RWL1$RBL1);
    if (WBL==1'b0 && WWL==1'b0 && RWL1==1'b0 )
       (RWL2 *> RBL2) = (tplh$RWL2$RBL2, tphl$RWL2$RBL2, tpxh$RWL2$RBL2, tphx$RWL2$RBL2, tplx$RWL2$RBL2, tpxl$RWL2$RBL2);
    if (WBL==1'b0 && WWL==1'b0 && RWL2==1'b1 )
       (RWL1 *> RBL1) = (tplh$RWL1$RBL1, tphl$RWL1$RBL1, tpxh$RWL1$RBL1, tphx$RWL1$RBL1, tplx$RWL1$RBL1, tpxl$RWL1$RBL1);
    if (WBL==1'b0 && WWL==1'b0 && RWL1==1'b1 )
       (RWL2 *> RBL2) = (tplh$RWL2$RBL2, tphl$RWL2$RBL2, tpxh$RWL2$RBL2, tphx$RWL2$RBL2, tplx$RWL2$RBL2, tpxl$RWL2$RBL2);
    if (WBL==1'b1 && WWL==1'b0 && RWL2==1'b0 )
       (RWL1 *> RBL1) = (tplh$RWL1$RBL1, tphl$RWL1$RBL1, tpxh$RWL1$RBL1, tphx$RWL1$RBL1, tplx$RWL1$RBL1, tpxl$RWL1$RBL1);
    if (WBL==1'b1 && WWL==1'b0 && RWL1==1'b0 )
       (RWL2 *> RBL2) = (tplh$RWL2$RBL2, tphl$RWL2$RBL2, tpxh$RWL2$RBL2, tphx$RWL2$RBL2, tplx$RWL2$RBL2, tpxl$RWL2$RBL2);
    if (WBL==1'b1 && WWL==1'b0 && RWL2==1'b1 )
       (RWL1 *> RBL1) = (tplh$RWL1$RBL1, tphl$RWL1$RBL1, tpxh$RWL1$RBL1, tphx$RWL1$RBL1, tplx$RWL1$RBL1, tpxl$RWL1$RBL1);
    if (WBL==1'b1 && WWL==1'b0 && RWL1==1'b1 )
       (RWL2 *> RBL2) = (tplh$RWL2$RBL2, tphl$RWL2$RBL2, tpxh$RWL2$RBL2, tphx$RWL2$RBL2, tplx$RWL2$RBL2, tpxl$RWL2$RBL2);
    if (WWL==1'b1 && RWL2==1'b0 )
       (RWL1 *> RBL1) = (tplh$RWL1$RBL1, tphl$RWL1$RBL1, tpxh$RWL1$RBL1, tphx$RWL1$RBL1, tplx$RWL1$RBL1, tpxl$RWL1$RBL1);
    if (WWL==1'b1 && RWL1==1'b0 )
       (RWL2 *> RBL2) = (tplh$RWL2$RBL2, tphl$RWL2$RBL2, tpxh$RWL2$RBL2, tphx$RWL2$RBL2, tplx$RWL2$RBL2, tpxl$RWL2$RBL2);
    if (WWL==1'b1 &&  RWL2==1'b0 )
       (WBL *> RBL1) = (tplh$WBL$RBL1, tphl$WBL$RBL1);
    if (WWL==1'b1 && RWL1==1'b0 )
       (WBL *> RBL2) = (tplh$WBL$RBL2, tphl$WBL$RBL2);
    if (WWL==1'b1 && RWL2==1'b1 )
       (RWL1 *> RBL1) = (tplh$RWL1$RBL1, tphl$RWL1$RBL1, tpxh$RWL1$RBL1, tphx$RWL1$RBL1, tplx$RWL1$RBL1, tpxl$RWL1$RBL1);
    if (WWL==1'b1 && RWL1==1'b1 )
       (RWL2 *> RBL2) = (tplh$RWL2$RBL2, tphl$RWL2$RBL2, tpxh$RWL2$RBL2, tphx$RWL2$RBL2, tplx$RWL2$RBL2, tpxl$RWL2$RBL2);
    if (WWL==1'b1 &&  RWL2==1'b1 )
       (WBL *> RBL1) = (tplh$WBL$RBL1, tphl$WBL$RBL1);
    if (WWL==1'b1 && RWL1==1'b1 )
       (WBL *> RBL2) = (tplh$WBL$RBL2, tphl$WBL$RBL2);
 

  endspecify

endmodule // RF2R1WSX1P4MA10TR
`endcelldefine
//$Id: rf.genpp,v 1.11 2006/05/18 09:44:11 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module RF2R1WSX1MA10TR (RBL1, RBL2, WBL, WWL, RWL1, RWL2);
output RBL1, RBL2;
input WBL, WWL, RWL1, RWL2;
reg NOTIFIER;

   not        I0 (WWLN, WWL);
   not        I1 (R1WN, RWL1);
   not        I2 (RWL2N, RWL2);
   udp_tlatrf I3 (n0, WBL, WWL, WWLN, NOTIFIER);
   bufif1     I4 (RBL1, n0, n2);
   bufif1     I5 (RBL2, n0, n3);
   udp_outrf  I6 (n2, n0, R1WN, RWL1);
   udp_outrf  I7 (n3, n0, RWL2N, RWL2);

  specify
    // delay parameters
    specparam
      tplh$WBL$RBL1 = 1.0,
      tphl$WBL$RBL1 = 1.0,
      tpxh$WBL$RBL1 = 1.0,
      tphx$WBL$RBL1 = 1.0,
      tplx$WBL$RBL1 = 1.0,
      tpxl$WBL$RBL1 = 1.0,
      tplh$WWL$RBL1 = 1.0,
      tphl$WWL$RBL1 = 1.0,
      tpxh$WWL$RBL1 = 1.0,
      tphx$WWL$RBL1 = 1.0,
      tplx$WWL$RBL1 = 1.0,
      tpxl$WWL$RBL1 = 1.0,
      tplh$RWL1$RBL1 = 1.0,
      tphl$RWL1$RBL1 = 1.0,
      tpxh$RWL1$RBL1 = 1.0,
      tphx$RWL1$RBL1 = 1.0,
      tplx$RWL1$RBL1 = 1.0,
      tpxl$RWL1$RBL1 = 1.0,
      tplh$RWL2$RBL1 = 1.0,
      tphl$RWL2$RBL1 = 1.0,
      tpxh$RWL2$RBL1 = 1.0,
      tphx$RWL2$RBL1 = 1.0,
      tplx$RWL2$RBL1 = 1.0,
      tpxl$RWL2$RBL1 = 1.0,
      tplh$WBL$RBL2 = 1.0,
      tphl$WBL$RBL2 = 1.0,
      tpxh$WBL$RBL2 = 1.0,
      tphx$WBL$RBL2 = 1.0,
      tplx$WBL$RBL2 = 1.0,
      tpxl$WBL$RBL2 = 1.0,
      tplh$WWL$RBL2 = 1.0,
      tphl$WWL$RBL2 = 1.0,
      tpxh$WWL$RBL2 = 1.0,
      tphx$WWL$RBL2 = 1.0,
      tplx$WWL$RBL2 = 1.0,
      tpxl$WWL$RBL2 = 1.0,
      tplh$RWL1$RBL2 = 1.0,
      tphl$RWL1$RBL2 = 1.0,
      tpxh$RWL1$RBL2 = 1.0,
      tphx$RWL1$RBL2 = 1.0,
      tplx$RWL1$RBL2 = 1.0,
      tpxl$RWL1$RBL2 = 1.0,
      tplh$RWL2$RBL2 = 1.0,
      tphl$RWL2$RBL2 = 1.0,
      tpxh$RWL2$RBL2 = 1.0,
      tphx$RWL2$RBL2 = 1.0,
      tplx$RWL2$RBL2 = 1.0,
      tpxl$RWL2$RBL2 = 1.0,
    tminpwh$WWL    = 1.0,
    tperiod$WWL    = 1.0,
    tsetup$WWL$WBL = 1.0,
    thold$WWL$WBL  = 0.5;

      // path delays
      ( WWL *> RBL1) = (tplh$WWL$RBL1, tphl$WWL$RBL1);
      ( WWL *> RBL2) = (tplh$WWL$RBL2, tphl$WWL$RBL2);
 
      // timing checks
      $width(posedge WWL, tminpwh$WWL, 0, NOTIFIER);
      $period(posedge WWL, tperiod$WWL, NOTIFIER);
      $setuphold(negedge WWL, posedge WBL, tsetup$WWL$WBL, thold$WWL$WBL, NOTIFIER);
      $setuphold(negedge WWL, negedge WBL, tsetup$WWL$WBL, thold$WWL$WBL, NOTIFIER);
    if (WBL==1'b0 && WWL==1'b0 && RWL2==1'b0 )
       (RWL1 *> RBL1) = (tplh$RWL1$RBL1, tphl$RWL1$RBL1, tpxh$RWL1$RBL1, tphx$RWL1$RBL1, tplx$RWL1$RBL1, tpxl$RWL1$RBL1);
    if (WBL==1'b0 && WWL==1'b0 && RWL1==1'b0 )
       (RWL2 *> RBL2) = (tplh$RWL2$RBL2, tphl$RWL2$RBL2, tpxh$RWL2$RBL2, tphx$RWL2$RBL2, tplx$RWL2$RBL2, tpxl$RWL2$RBL2);
    if (WBL==1'b0 && WWL==1'b0 && RWL2==1'b1 )
       (RWL1 *> RBL1) = (tplh$RWL1$RBL1, tphl$RWL1$RBL1, tpxh$RWL1$RBL1, tphx$RWL1$RBL1, tplx$RWL1$RBL1, tpxl$RWL1$RBL1);
    if (WBL==1'b0 && WWL==1'b0 && RWL1==1'b1 )
       (RWL2 *> RBL2) = (tplh$RWL2$RBL2, tphl$RWL2$RBL2, tpxh$RWL2$RBL2, tphx$RWL2$RBL2, tplx$RWL2$RBL2, tpxl$RWL2$RBL2);
    if (WBL==1'b1 && WWL==1'b0 && RWL2==1'b0 )
       (RWL1 *> RBL1) = (tplh$RWL1$RBL1, tphl$RWL1$RBL1, tpxh$RWL1$RBL1, tphx$RWL1$RBL1, tplx$RWL1$RBL1, tpxl$RWL1$RBL1);
    if (WBL==1'b1 && WWL==1'b0 && RWL1==1'b0 )
       (RWL2 *> RBL2) = (tplh$RWL2$RBL2, tphl$RWL2$RBL2, tpxh$RWL2$RBL2, tphx$RWL2$RBL2, tplx$RWL2$RBL2, tpxl$RWL2$RBL2);
    if (WBL==1'b1 && WWL==1'b0 && RWL2==1'b1 )
       (RWL1 *> RBL1) = (tplh$RWL1$RBL1, tphl$RWL1$RBL1, tpxh$RWL1$RBL1, tphx$RWL1$RBL1, tplx$RWL1$RBL1, tpxl$RWL1$RBL1);
    if (WBL==1'b1 && WWL==1'b0 && RWL1==1'b1 )
       (RWL2 *> RBL2) = (tplh$RWL2$RBL2, tphl$RWL2$RBL2, tpxh$RWL2$RBL2, tphx$RWL2$RBL2, tplx$RWL2$RBL2, tpxl$RWL2$RBL2);
    if (WWL==1'b1 && RWL2==1'b0 )
       (RWL1 *> RBL1) = (tplh$RWL1$RBL1, tphl$RWL1$RBL1, tpxh$RWL1$RBL1, tphx$RWL1$RBL1, tplx$RWL1$RBL1, tpxl$RWL1$RBL1);
    if (WWL==1'b1 && RWL1==1'b0 )
       (RWL2 *> RBL2) = (tplh$RWL2$RBL2, tphl$RWL2$RBL2, tpxh$RWL2$RBL2, tphx$RWL2$RBL2, tplx$RWL2$RBL2, tpxl$RWL2$RBL2);
    if (WWL==1'b1 &&  RWL2==1'b0 )
       (WBL *> RBL1) = (tplh$WBL$RBL1, tphl$WBL$RBL1);
    if (WWL==1'b1 && RWL1==1'b0 )
       (WBL *> RBL2) = (tplh$WBL$RBL2, tphl$WBL$RBL2);
    if (WWL==1'b1 && RWL2==1'b1 )
       (RWL1 *> RBL1) = (tplh$RWL1$RBL1, tphl$RWL1$RBL1, tpxh$RWL1$RBL1, tphx$RWL1$RBL1, tplx$RWL1$RBL1, tpxl$RWL1$RBL1);
    if (WWL==1'b1 && RWL1==1'b1 )
       (RWL2 *> RBL2) = (tplh$RWL2$RBL2, tphl$RWL2$RBL2, tpxh$RWL2$RBL2, tphx$RWL2$RBL2, tplx$RWL2$RBL2, tpxl$RWL2$RBL2);
    if (WWL==1'b1 &&  RWL2==1'b1 )
       (WBL *> RBL1) = (tplh$WBL$RBL1, tphl$WBL$RBL1);
    if (WWL==1'b1 && RWL1==1'b1 )
       (WBL *> RBL2) = (tplh$WBL$RBL2, tphl$WBL$RBL2);
 

  endspecify

endmodule // RF2R1WSX1MA10TR
`endcelldefine
//$Id: rf.genpp,v 1.11 2006/05/18 09:44:11 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module RF1R2WSX2MA10TR (RBL, WBL1, WWL1, WBL2, WWL2, RWL);
output RBL;
input WBL1, WWL1, WBL2, WWL2, RWL;
reg NOTIFIER;

   not I0 (ckn, ck);
   or  I1 (ck, WWL1, WWL2); 
   udp_wao I2 (wr, WBL1, WBL2, WWL1, WWL2);
   udp_tlatrf I3 (n0, wr, ck, ckn, NOTIFIER);
   not I4 (n1, n0);
   notif1 I5 (RBL, n1, RWL);

  specify
    // delay parameters
    specparam
      tplh$WBL1$RBL = 1.0,
      tphl$WBL1$RBL = 1.0,
      tpxh$WBL1$RBL = 1.0,
      tphx$WBL1$RBL = 1.0,
      tplx$WBL1$RBL = 1.0,
      tpxl$WBL1$RBL = 1.0,
      tplh$WWL1$RBL = 1.0,
      tphl$WWL1$RBL = 1.0,
      tpxh$WWL1$RBL = 1.0,
      tphx$WWL1$RBL = 1.0,
      tplx$WWL1$RBL = 1.0,
      tpxl$WWL1$RBL = 1.0,
      tplh$WBL2$RBL = 1.0,
      tphl$WBL2$RBL = 1.0,
      tpxh$WBL2$RBL = 1.0,
      tphx$WBL2$RBL = 1.0,
      tplx$WBL2$RBL = 1.0,
      tpxl$WBL2$RBL = 1.0,
      tplh$WWL2$RBL = 1.0,
      tphl$WWL2$RBL = 1.0,
      tpxh$WWL2$RBL = 1.0,
      tphx$WWL2$RBL = 1.0,
      tplx$WWL2$RBL = 1.0,
      tpxl$WWL2$RBL = 1.0,
      tplh$RWL$RBL = 1.0,
      tphl$RWL$RBL = 1.0,
      tpxh$RWL$RBL = 1.0,
      tphx$RWL$RBL = 1.0,
      tplx$RWL$RBL = 1.0,
      tpxl$RWL$RBL = 1.0,
    tsetup$WWL1$WBL1 = 1.0,
    thold$WWL1$WBL1  = 0.5,
    tsetup$WWL2$WBL2 = 1.0,
    thold$WWL2$WBL2  = 0.5,
    tminpwh$WWL1    = 1.0,
    tperiod$WWL1    = 1.0,
    tminpwh$WWL2    = 1.0,
    tperiod$WWL2    = 1.0;

      // path delays
 
      // timing checks
      $setuphold(negedge WWL1, posedge WBL1, tsetup$WWL1$WBL1, thold$WWL1$WBL1, NOTIFIER);
      $setuphold(negedge WWL1, negedge WBL1, tsetup$WWL1$WBL1, thold$WWL1$WBL1, NOTIFIER);
      $setuphold(negedge WWL2, posedge WBL2, tsetup$WWL2$WBL2, thold$WWL2$WBL2, NOTIFIER);
      $setuphold(negedge WWL2, negedge WBL2, tsetup$WWL2$WBL2, thold$WWL2$WBL2, NOTIFIER);
      $width(posedge WWL1, tminpwh$WWL1, 0, NOTIFIER);
      $period(posedge WWL1, tperiod$WWL1, NOTIFIER);
      $width(posedge WWL2, tminpwh$WWL2, 0, NOTIFIER);
      $period(posedge WWL2, tperiod$WWL2, NOTIFIER);
    if (WWL2 == 1'b0 && RWL == 1'b1 )
       (posedge  WWL1 *> (RBL -: WBL1)) = (tplh$WWL1$RBL, tphl$WWL1$RBL);
    if (WWL1 == 1'b0 && RWL == 1'b1 )
       (posedge  WWL2 *> (RBL -: WBL2)) = (tplh$WWL2$RBL, tphl$WWL2$RBL);
    if (WWL1 == 1'b1 && WWL2 == 1'b0 && RWL == 1'b1 )
       (WBL1 *> RBL) = (tplh$WBL1$RBL, tphl$WBL1$RBL);
    if (WWL1 == 1'b0 && WWL2 == 1'b1 && RWL == 1'b1 )
       (WBL2 *> RBL) = (tplh$WBL2$RBL, tphl$WBL2$RBL);
    if (WWL1 == 1'b0 && WWL2 == 1'b0 )
       (RWL *> RBL) = (tplh$RWL$RBL, tphl$RWL$RBL, tpxh$RWL$RBL, tphx$RWL$RBL, tplx$RWL$RBL, tpxl$RWL$RBL);
    if (WWL1 == 1'b0 && WWL2 == 1'b1 )
       (RWL *> RBL) = (tplh$RWL$RBL, tphl$RWL$RBL, tpxh$RWL$RBL, tphx$RWL$RBL, tplx$RWL$RBL, tpxl$RWL$RBL);
    if (WWL1 == 1'b1 && WWL2 == 1'b0 )
       (RWL *> RBL) = (tplh$RWL$RBL, tphl$RWL$RBL, tpxh$RWL$RBL, tphx$RWL$RBL, tplx$RWL$RBL, tpxl$RWL$RBL);
    if (WWL1 == 1'b1 && WWL2 == 1'b1 )
       (RWL *> RBL) = (tplh$RWL$RBL, tphl$RWL$RBL, tpxh$RWL$RBL, tphx$RWL$RBL, tplx$RWL$RBL, tpxl$RWL$RBL);
 

  endspecify

endmodule // RF1R2WSX2MA10TR
`endcelldefine
//$Id: rf.genpp,v 1.11 2006/05/18 09:44:11 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module RF1R2WSX1P4MA10TR (RBL, WBL1, WWL1, WBL2, WWL2, RWL);
output RBL;
input WBL1, WWL1, WBL2, WWL2, RWL;
reg NOTIFIER;

   not I0 (ckn, ck);
   or  I1 (ck, WWL1, WWL2); 
   udp_wao I2 (wr, WBL1, WBL2, WWL1, WWL2);
   udp_tlatrf I3 (n0, wr, ck, ckn, NOTIFIER);
   not I4 (n1, n0);
   notif1 I5 (RBL, n1, RWL);

  specify
    // delay parameters
    specparam
      tplh$WBL1$RBL = 1.0,
      tphl$WBL1$RBL = 1.0,
      tpxh$WBL1$RBL = 1.0,
      tphx$WBL1$RBL = 1.0,
      tplx$WBL1$RBL = 1.0,
      tpxl$WBL1$RBL = 1.0,
      tplh$WWL1$RBL = 1.0,
      tphl$WWL1$RBL = 1.0,
      tpxh$WWL1$RBL = 1.0,
      tphx$WWL1$RBL = 1.0,
      tplx$WWL1$RBL = 1.0,
      tpxl$WWL1$RBL = 1.0,
      tplh$WBL2$RBL = 1.0,
      tphl$WBL2$RBL = 1.0,
      tpxh$WBL2$RBL = 1.0,
      tphx$WBL2$RBL = 1.0,
      tplx$WBL2$RBL = 1.0,
      tpxl$WBL2$RBL = 1.0,
      tplh$WWL2$RBL = 1.0,
      tphl$WWL2$RBL = 1.0,
      tpxh$WWL2$RBL = 1.0,
      tphx$WWL2$RBL = 1.0,
      tplx$WWL2$RBL = 1.0,
      tpxl$WWL2$RBL = 1.0,
      tplh$RWL$RBL = 1.0,
      tphl$RWL$RBL = 1.0,
      tpxh$RWL$RBL = 1.0,
      tphx$RWL$RBL = 1.0,
      tplx$RWL$RBL = 1.0,
      tpxl$RWL$RBL = 1.0,
    tsetup$WWL1$WBL1 = 1.0,
    thold$WWL1$WBL1  = 0.5,
    tsetup$WWL2$WBL2 = 1.0,
    thold$WWL2$WBL2  = 0.5,
    tminpwh$WWL1    = 1.0,
    tperiod$WWL1    = 1.0,
    tminpwh$WWL2    = 1.0,
    tperiod$WWL2    = 1.0;

      // path delays
 
      // timing checks
      $setuphold(negedge WWL1, posedge WBL1, tsetup$WWL1$WBL1, thold$WWL1$WBL1, NOTIFIER);
      $setuphold(negedge WWL1, negedge WBL1, tsetup$WWL1$WBL1, thold$WWL1$WBL1, NOTIFIER);
      $setuphold(negedge WWL2, posedge WBL2, tsetup$WWL2$WBL2, thold$WWL2$WBL2, NOTIFIER);
      $setuphold(negedge WWL2, negedge WBL2, tsetup$WWL2$WBL2, thold$WWL2$WBL2, NOTIFIER);
      $width(posedge WWL1, tminpwh$WWL1, 0, NOTIFIER);
      $period(posedge WWL1, tperiod$WWL1, NOTIFIER);
      $width(posedge WWL2, tminpwh$WWL2, 0, NOTIFIER);
      $period(posedge WWL2, tperiod$WWL2, NOTIFIER);
    if (WWL2 == 1'b0 && RWL == 1'b1 )
       (posedge  WWL1 *> (RBL -: WBL1)) = (tplh$WWL1$RBL, tphl$WWL1$RBL);
    if (WWL1 == 1'b0 && RWL == 1'b1 )
       (posedge  WWL2 *> (RBL -: WBL2)) = (tplh$WWL2$RBL, tphl$WWL2$RBL);
    if (WWL1 == 1'b1 && WWL2 == 1'b0 && RWL == 1'b1 )
       (WBL1 *> RBL) = (tplh$WBL1$RBL, tphl$WBL1$RBL);
    if (WWL1 == 1'b0 && WWL2 == 1'b1 && RWL == 1'b1 )
       (WBL2 *> RBL) = (tplh$WBL2$RBL, tphl$WBL2$RBL);
    if (WWL1 == 1'b0 && WWL2 == 1'b0 )
       (RWL *> RBL) = (tplh$RWL$RBL, tphl$RWL$RBL, tpxh$RWL$RBL, tphx$RWL$RBL, tplx$RWL$RBL, tpxl$RWL$RBL);
    if (WWL1 == 1'b0 && WWL2 == 1'b1 )
       (RWL *> RBL) = (tplh$RWL$RBL, tphl$RWL$RBL, tpxh$RWL$RBL, tphx$RWL$RBL, tplx$RWL$RBL, tpxl$RWL$RBL);
    if (WWL1 == 1'b1 && WWL2 == 1'b0 )
       (RWL *> RBL) = (tplh$RWL$RBL, tphl$RWL$RBL, tpxh$RWL$RBL, tphx$RWL$RBL, tplx$RWL$RBL, tpxl$RWL$RBL);
    if (WWL1 == 1'b1 && WWL2 == 1'b1 )
       (RWL *> RBL) = (tplh$RWL$RBL, tphl$RWL$RBL, tpxh$RWL$RBL, tphx$RWL$RBL, tplx$RWL$RBL, tpxl$RWL$RBL);
 

  endspecify

endmodule // RF1R2WSX1P4MA10TR
`endcelldefine
//$Id: rf.genpp,v 1.11 2006/05/18 09:44:11 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module RF1R2WSX1MA10TR (RBL, WBL1, WWL1, WBL2, WWL2, RWL);
output RBL;
input WBL1, WWL1, WBL2, WWL2, RWL;
reg NOTIFIER;

   not I0 (ckn, ck);
   or  I1 (ck, WWL1, WWL2); 
   udp_wao I2 (wr, WBL1, WBL2, WWL1, WWL2);
   udp_tlatrf I3 (n0, wr, ck, ckn, NOTIFIER);
   not I4 (n1, n0);
   notif1 I5 (RBL, n1, RWL);

  specify
    // delay parameters
    specparam
      tplh$WBL1$RBL = 1.0,
      tphl$WBL1$RBL = 1.0,
      tpxh$WBL1$RBL = 1.0,
      tphx$WBL1$RBL = 1.0,
      tplx$WBL1$RBL = 1.0,
      tpxl$WBL1$RBL = 1.0,
      tplh$WWL1$RBL = 1.0,
      tphl$WWL1$RBL = 1.0,
      tpxh$WWL1$RBL = 1.0,
      tphx$WWL1$RBL = 1.0,
      tplx$WWL1$RBL = 1.0,
      tpxl$WWL1$RBL = 1.0,
      tplh$WBL2$RBL = 1.0,
      tphl$WBL2$RBL = 1.0,
      tpxh$WBL2$RBL = 1.0,
      tphx$WBL2$RBL = 1.0,
      tplx$WBL2$RBL = 1.0,
      tpxl$WBL2$RBL = 1.0,
      tplh$WWL2$RBL = 1.0,
      tphl$WWL2$RBL = 1.0,
      tpxh$WWL2$RBL = 1.0,
      tphx$WWL2$RBL = 1.0,
      tplx$WWL2$RBL = 1.0,
      tpxl$WWL2$RBL = 1.0,
      tplh$RWL$RBL = 1.0,
      tphl$RWL$RBL = 1.0,
      tpxh$RWL$RBL = 1.0,
      tphx$RWL$RBL = 1.0,
      tplx$RWL$RBL = 1.0,
      tpxl$RWL$RBL = 1.0,
    tsetup$WWL1$WBL1 = 1.0,
    thold$WWL1$WBL1  = 0.5,
    tsetup$WWL2$WBL2 = 1.0,
    thold$WWL2$WBL2  = 0.5,
    tminpwh$WWL1    = 1.0,
    tperiod$WWL1    = 1.0,
    tminpwh$WWL2    = 1.0,
    tperiod$WWL2    = 1.0;

      // path delays
 
      // timing checks
      $setuphold(negedge WWL1, posedge WBL1, tsetup$WWL1$WBL1, thold$WWL1$WBL1, NOTIFIER);
      $setuphold(negedge WWL1, negedge WBL1, tsetup$WWL1$WBL1, thold$WWL1$WBL1, NOTIFIER);
      $setuphold(negedge WWL2, posedge WBL2, tsetup$WWL2$WBL2, thold$WWL2$WBL2, NOTIFIER);
      $setuphold(negedge WWL2, negedge WBL2, tsetup$WWL2$WBL2, thold$WWL2$WBL2, NOTIFIER);
      $width(posedge WWL1, tminpwh$WWL1, 0, NOTIFIER);
      $period(posedge WWL1, tperiod$WWL1, NOTIFIER);
      $width(posedge WWL2, tminpwh$WWL2, 0, NOTIFIER);
      $period(posedge WWL2, tperiod$WWL2, NOTIFIER);
    if (WWL2 == 1'b0 && RWL == 1'b1 )
       (posedge  WWL1 *> (RBL -: WBL1)) = (tplh$WWL1$RBL, tphl$WWL1$RBL);
    if (WWL1 == 1'b0 && RWL == 1'b1 )
       (posedge  WWL2 *> (RBL -: WBL2)) = (tplh$WWL2$RBL, tphl$WWL2$RBL);
    if (WWL1 == 1'b1 && WWL2 == 1'b0 && RWL == 1'b1 )
       (WBL1 *> RBL) = (tplh$WBL1$RBL, tphl$WBL1$RBL);
    if (WWL1 == 1'b0 && WWL2 == 1'b1 && RWL == 1'b1 )
       (WBL2 *> RBL) = (tplh$WBL2$RBL, tphl$WBL2$RBL);
    if (WWL1 == 1'b0 && WWL2 == 1'b0 )
       (RWL *> RBL) = (tplh$RWL$RBL, tphl$RWL$RBL, tpxh$RWL$RBL, tphx$RWL$RBL, tplx$RWL$RBL, tpxl$RWL$RBL);
    if (WWL1 == 1'b0 && WWL2 == 1'b1 )
       (RWL *> RBL) = (tplh$RWL$RBL, tphl$RWL$RBL, tpxh$RWL$RBL, tphx$RWL$RBL, tplx$RWL$RBL, tpxl$RWL$RBL);
    if (WWL1 == 1'b1 && WWL2 == 1'b0 )
       (RWL *> RBL) = (tplh$RWL$RBL, tphl$RWL$RBL, tpxh$RWL$RBL, tphx$RWL$RBL, tplx$RWL$RBL, tpxl$RWL$RBL);
    if (WWL1 == 1'b1 && WWL2 == 1'b1 )
       (RWL *> RBL) = (tplh$RWL$RBL, tphl$RWL$RBL, tpxh$RWL$RBL, tphx$RWL$RBL, tplx$RWL$RBL, tpxl$RWL$RBL);
 

  endspecify

endmodule // RF1R2WSX1MA10TR
`endcelldefine
//$Id: rf.genpp,v 1.11 2006/05/18 09:44:11 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module RF1R1WSX2MA10TR (RBL, WBL, WWL, RWL);
output RBL;
input WBL, WWL, RWL;
reg NOTIFIER;

   not II (wwn,WWL);
   udp_tlatrf I0 (n0, WBL, WWL, wwn, NOTIFIER);
   bufif1     I1 (RBL, n0, RWL);

  specify
    // delay parameters
    specparam
      tplh$WBL$RBL = 1.0,
      tphl$WBL$RBL = 1.0,
      tplh$WWL$RBL = 1.0,
      tphl$WWL$RBL = 1.0,
      tplh$RWL$RBL = 1.0,
      tphl$RWL$RBL = 1.0,
    tsetup$WWL$WBL = 1.0,
    thold$WWL$WBL  = 0.5,
    tminpwh$WWL    = 1.0,
    tperiod$WWL    = 1.0;

      // path delays
      ( posedge WWL *> (RBL -:WBL )) = (tplh$WWL$RBL, tphl$WWL$RBL);
      ( WBL *> RBL ) = (tplh$WBL$RBL, tphl$WBL$RBL);
      ( RWL *> RBL ) = (tplh$RWL$RBL, tphl$RWL$RBL);
 
      // timing checks
      $width(posedge WWL, tminpwh$WWL, 0, NOTIFIER);
      $period(posedge WWL, tperiod$WWL, NOTIFIER);
      $setuphold(negedge WWL, posedge WBL, tsetup$WWL$WBL, thold$WWL$WBL, NOTIFIER);
      $setuphold(negedge WWL, negedge WBL, tsetup$WWL$WBL, thold$WWL$WBL, NOTIFIER);
 

  endspecify

endmodule // RF1R1WSX2MA10TR
`endcelldefine
//$Id: rf.genpp,v 1.11 2006/05/18 09:44:11 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module RF1R1WSX1P4MA10TR (RBL, WBL, WWL, RWL);
output RBL;
input WBL, WWL, RWL;
reg NOTIFIER;

   not II (wwn,WWL);
   udp_tlatrf I0 (n0, WBL, WWL, wwn, NOTIFIER);
   bufif1     I1 (RBL, n0, RWL);

  specify
    // delay parameters
    specparam
      tplh$WBL$RBL = 1.0,
      tphl$WBL$RBL = 1.0,
      tplh$WWL$RBL = 1.0,
      tphl$WWL$RBL = 1.0,
      tplh$RWL$RBL = 1.0,
      tphl$RWL$RBL = 1.0,
    tsetup$WWL$WBL = 1.0,
    thold$WWL$WBL  = 0.5,
    tminpwh$WWL    = 1.0,
    tperiod$WWL    = 1.0;

      // path delays
      ( posedge WWL *> (RBL -:WBL )) = (tplh$WWL$RBL, tphl$WWL$RBL);
      ( WBL *> RBL ) = (tplh$WBL$RBL, tphl$WBL$RBL);
      ( RWL *> RBL ) = (tplh$RWL$RBL, tphl$RWL$RBL);
 
      // timing checks
      $width(posedge WWL, tminpwh$WWL, 0, NOTIFIER);
      $period(posedge WWL, tperiod$WWL, NOTIFIER);
      $setuphold(negedge WWL, posedge WBL, tsetup$WWL$WBL, thold$WWL$WBL, NOTIFIER);
      $setuphold(negedge WWL, negedge WBL, tsetup$WWL$WBL, thold$WWL$WBL, NOTIFIER);
 

  endspecify

endmodule // RF1R1WSX1P4MA10TR
`endcelldefine
//$Id: rf.genpp,v 1.11 2006/05/18 09:44:11 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module RF1R1WSX1MA10TR (RBL, WBL, WWL, RWL);
output RBL;
input WBL, WWL, RWL;
reg NOTIFIER;

   not II (wwn,WWL);
   udp_tlatrf I0 (n0, WBL, WWL, wwn, NOTIFIER);
   bufif1     I1 (RBL, n0, RWL);

  specify
    // delay parameters
    specparam
      tplh$WBL$RBL = 1.0,
      tphl$WBL$RBL = 1.0,
      tplh$WWL$RBL = 1.0,
      tphl$WWL$RBL = 1.0,
      tplh$RWL$RBL = 1.0,
      tphl$RWL$RBL = 1.0,
    tsetup$WWL$WBL = 1.0,
    thold$WWL$WBL  = 0.5,
    tminpwh$WWL    = 1.0,
    tperiod$WWL    = 1.0;

      // path delays
      ( posedge WWL *> (RBL -:WBL )) = (tplh$WWL$RBL, tphl$WWL$RBL);
      ( WBL *> RBL ) = (tplh$WBL$RBL, tphl$WBL$RBL);
      ( RWL *> RBL ) = (tplh$RWL$RBL, tphl$RWL$RBL);
 
      // timing checks
      $width(posedge WWL, tminpwh$WWL, 0, NOTIFIER);
      $period(posedge WWL, tperiod$WWL, NOTIFIER);
      $setuphold(negedge WWL, posedge WBL, tsetup$WWL$WBL, thold$WWL$WBL, NOTIFIER);
      $setuphold(negedge WWL, negedge WBL, tsetup$WWL$WBL, thold$WWL$WBL, NOTIFIER);
 

  endspecify

endmodule // RF1R1WSX1MA10TR
`endcelldefine
//$Id: ckgate.genpp,v 1.15 2006/06/21 06:18:22 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module PREICGX9BA10TR (ECK, E, SE, CK);
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, NOTIFIER);
  and      I2 (ECK, n0, CK);
  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SE$ECK   = 1.0,
      tphl$SE$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SE$CK  = 1.0,
      thold$SE$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      if (E==1'b0 && SE==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b0 && SE==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SE==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SE==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SE == 0), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (SE == 0), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
    $setuphold(posedge CK, posedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER);
    $setuphold(posedge CK, negedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER);
  endspecify

endmodule //PREICGX9BA10TR
`endcelldefine
//$Id: ckgate.genpp,v 1.15 2006/06/21 06:18:22 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module PREICGX7P5BA10TR (ECK, E, SE, CK);
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, NOTIFIER);
  and      I2 (ECK, n0, CK);
  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SE$ECK   = 1.0,
      tphl$SE$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SE$CK  = 1.0,
      thold$SE$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      if (E==1'b0 && SE==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b0 && SE==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SE==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SE==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SE == 0), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (SE == 0), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
    $setuphold(posedge CK, posedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER);
    $setuphold(posedge CK, negedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER);
  endspecify

endmodule //PREICGX7P5BA10TR
`endcelldefine
//$Id: ckgate.genpp,v 1.15 2006/06/21 06:18:22 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module PREICGX6BA10TR (ECK, E, SE, CK);
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, NOTIFIER);
  and      I2 (ECK, n0, CK);
  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SE$ECK   = 1.0,
      tphl$SE$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SE$CK  = 1.0,
      thold$SE$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      if (E==1'b0 && SE==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b0 && SE==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SE==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SE==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SE == 0), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (SE == 0), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
    $setuphold(posedge CK, posedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER);
    $setuphold(posedge CK, negedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER);
  endspecify

endmodule //PREICGX6BA10TR
`endcelldefine
//$Id: ckgate.genpp,v 1.15 2006/06/21 06:18:22 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module PREICGX5BA10TR (ECK, E, SE, CK);
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, NOTIFIER);
  and      I2 (ECK, n0, CK);
  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SE$ECK   = 1.0,
      tphl$SE$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SE$CK  = 1.0,
      thold$SE$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      if (E==1'b0 && SE==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b0 && SE==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SE==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SE==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SE == 0), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (SE == 0), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
    $setuphold(posedge CK, posedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER);
    $setuphold(posedge CK, negedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER);
  endspecify

endmodule //PREICGX5BA10TR
`endcelldefine
//$Id: ckgate.genpp,v 1.15 2006/06/21 06:18:22 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module PREICGX4BA10TR (ECK, E, SE, CK);
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, NOTIFIER);
  and      I2 (ECK, n0, CK);
  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SE$ECK   = 1.0,
      tphl$SE$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SE$CK  = 1.0,
      thold$SE$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      if (E==1'b0 && SE==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b0 && SE==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SE==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SE==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SE == 0), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (SE == 0), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
    $setuphold(posedge CK, posedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER);
    $setuphold(posedge CK, negedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER);
  endspecify

endmodule //PREICGX4BA10TR
`endcelldefine
//$Id: ckgate.genpp,v 1.15 2006/06/21 06:18:22 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module PREICGX3P5BA10TR (ECK, E, SE, CK);
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, NOTIFIER);
  and      I2 (ECK, n0, CK);
  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SE$ECK   = 1.0,
      tphl$SE$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SE$CK  = 1.0,
      thold$SE$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      if (E==1'b0 && SE==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b0 && SE==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SE==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SE==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SE == 0), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (SE == 0), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
    $setuphold(posedge CK, posedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER);
    $setuphold(posedge CK, negedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER);
  endspecify

endmodule //PREICGX3P5BA10TR
`endcelldefine
//$Id: ckgate.genpp,v 1.15 2006/06/21 06:18:22 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module PREICGX3BA10TR (ECK, E, SE, CK);
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, NOTIFIER);
  and      I2 (ECK, n0, CK);
  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SE$ECK   = 1.0,
      tphl$SE$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SE$CK  = 1.0,
      thold$SE$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      if (E==1'b0 && SE==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b0 && SE==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SE==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SE==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SE == 0), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (SE == 0), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
    $setuphold(posedge CK, posedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER);
    $setuphold(posedge CK, negedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER);
  endspecify

endmodule //PREICGX3BA10TR
`endcelldefine
//$Id: ckgate.genpp,v 1.15 2006/06/21 06:18:22 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module PREICGX2P5BA10TR (ECK, E, SE, CK);
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, NOTIFIER);
  and      I2 (ECK, n0, CK);
  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SE$ECK   = 1.0,
      tphl$SE$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SE$CK  = 1.0,
      thold$SE$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      if (E==1'b0 && SE==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b0 && SE==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SE==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SE==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SE == 0), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (SE == 0), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
    $setuphold(posedge CK, posedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER);
    $setuphold(posedge CK, negedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER);
  endspecify

endmodule //PREICGX2P5BA10TR
`endcelldefine
//$Id: ckgate.genpp,v 1.15 2006/06/21 06:18:22 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module PREICGX2BA10TR (ECK, E, SE, CK);
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, NOTIFIER);
  and      I2 (ECK, n0, CK);
  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SE$ECK   = 1.0,
      tphl$SE$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SE$CK  = 1.0,
      thold$SE$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      if (E==1'b0 && SE==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b0 && SE==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SE==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SE==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SE == 0), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (SE == 0), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
    $setuphold(posedge CK, posedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER);
    $setuphold(posedge CK, negedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER);
  endspecify

endmodule //PREICGX2BA10TR
`endcelldefine
//$Id: ckgate.genpp,v 1.15 2006/06/21 06:18:22 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module PREICGX1P7BA10TR (ECK, E, SE, CK);
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, NOTIFIER);
  and      I2 (ECK, n0, CK);
  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SE$ECK   = 1.0,
      tphl$SE$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SE$CK  = 1.0,
      thold$SE$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      if (E==1'b0 && SE==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b0 && SE==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SE==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SE==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SE == 0), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (SE == 0), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
    $setuphold(posedge CK, posedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER);
    $setuphold(posedge CK, negedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER);
  endspecify

endmodule //PREICGX1P7BA10TR
`endcelldefine
//$Id: ckgate.genpp,v 1.15 2006/06/21 06:18:22 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module PREICGX1P4BA10TR (ECK, E, SE, CK);
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, NOTIFIER);
  and      I2 (ECK, n0, CK);
  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SE$ECK   = 1.0,
      tphl$SE$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SE$CK  = 1.0,
      thold$SE$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      if (E==1'b0 && SE==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b0 && SE==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SE==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SE==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SE == 0), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (SE == 0), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
    $setuphold(posedge CK, posedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER);
    $setuphold(posedge CK, negedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER);
  endspecify

endmodule //PREICGX1P4BA10TR
`endcelldefine
//$Id: ckgate.genpp,v 1.15 2006/06/21 06:18:22 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module PREICGX1P2BA10TR (ECK, E, SE, CK);
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, NOTIFIER);
  and      I2 (ECK, n0, CK);
  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SE$ECK   = 1.0,
      tphl$SE$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SE$CK  = 1.0,
      thold$SE$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      if (E==1'b0 && SE==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b0 && SE==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SE==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SE==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SE == 0), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (SE == 0), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
    $setuphold(posedge CK, posedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER);
    $setuphold(posedge CK, negedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER);
  endspecify

endmodule //PREICGX1P2BA10TR
`endcelldefine
//$Id: ckgate.genpp,v 1.15 2006/06/21 06:18:22 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module PREICGX1BA10TR (ECK, E, SE, CK);
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, NOTIFIER);
  and      I2 (ECK, n0, CK);
  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SE$ECK   = 1.0,
      tphl$SE$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SE$CK  = 1.0,
      thold$SE$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      if (E==1'b0 && SE==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b0 && SE==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SE==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SE==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SE == 0), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (SE == 0), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
    $setuphold(posedge CK, posedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER);
    $setuphold(posedge CK, negedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER);
  endspecify

endmodule //PREICGX1BA10TR
`endcelldefine
//$Id: ckgate.genpp,v 1.15 2006/06/21 06:18:22 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module PREICGX16BA10TR (ECK, E, SE, CK);
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, NOTIFIER);
  and      I2 (ECK, n0, CK);
  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SE$ECK   = 1.0,
      tphl$SE$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SE$CK  = 1.0,
      thold$SE$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      if (E==1'b0 && SE==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b0 && SE==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SE==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SE==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SE == 0), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (SE == 0), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
    $setuphold(posedge CK, posedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER);
    $setuphold(posedge CK, negedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER);
  endspecify

endmodule //PREICGX16BA10TR
`endcelldefine
//$Id: ckgate.genpp,v 1.15 2006/06/21 06:18:22 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module PREICGX13BA10TR (ECK, E, SE, CK);
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, NOTIFIER);
  and      I2 (ECK, n0, CK);
  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SE$ECK   = 1.0,
      tphl$SE$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SE$CK  = 1.0,
      thold$SE$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      if (E==1'b0 && SE==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b0 && SE==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SE==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SE==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SE == 0), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (SE == 0), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
    $setuphold(posedge CK, posedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER);
    $setuphold(posedge CK, negedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER);
  endspecify

endmodule //PREICGX13BA10TR
`endcelldefine
//$Id: ckgate.genpp,v 1.15 2006/06/21 06:18:22 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module PREICGX11BA10TR (ECK, E, SE, CK);
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, NOTIFIER);
  and      I2 (ECK, n0, CK);
  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SE$ECK   = 1.0,
      tphl$SE$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SE$CK  = 1.0,
      thold$SE$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      if (E==1'b0 && SE==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b0 && SE==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SE==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SE==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SE == 0), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (SE == 0), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
    $setuphold(posedge CK, posedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER);
    $setuphold(posedge CK, negedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER);
  endspecify

endmodule //PREICGX11BA10TR
`endcelldefine
//$Id: ckgate.genpp,v 1.15 2006/06/21 06:18:22 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module PREICGX0P8BA10TR (ECK, E, SE, CK);
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, NOTIFIER);
  and      I2 (ECK, n0, CK);
  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SE$ECK   = 1.0,
      tphl$SE$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SE$CK  = 1.0,
      thold$SE$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      if (E==1'b0 && SE==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b0 && SE==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SE==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SE==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SE == 0), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (SE == 0), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
    $setuphold(posedge CK, posedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER);
    $setuphold(posedge CK, negedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER);
  endspecify

endmodule //PREICGX0P8BA10TR
`endcelldefine
//$Id: ckgate.genpp,v 1.15 2006/06/21 06:18:22 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module PREICGX0P7BA10TR (ECK, E, SE, CK);
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, NOTIFIER);
  and      I2 (ECK, n0, CK);
  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SE$ECK   = 1.0,
      tphl$SE$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SE$CK  = 1.0,
      thold$SE$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      if (E==1'b0 && SE==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b0 && SE==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SE==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SE==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SE == 0), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (SE == 0), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
    $setuphold(posedge CK, posedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER);
    $setuphold(posedge CK, negedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER);
  endspecify

endmodule //PREICGX0P7BA10TR
`endcelldefine
//$Id: ckgate.genpp,v 1.15 2006/06/21 06:18:22 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module PREICGX0P6BA10TR (ECK, E, SE, CK);
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, NOTIFIER);
  and      I2 (ECK, n0, CK);
  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SE$ECK   = 1.0,
      tphl$SE$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SE$CK  = 1.0,
      thold$SE$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      if (E==1'b0 && SE==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b0 && SE==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SE==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SE==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SE == 0), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (SE == 0), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
    $setuphold(posedge CK, posedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER);
    $setuphold(posedge CK, negedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER);
  endspecify

endmodule //PREICGX0P6BA10TR
`endcelldefine
//$Id: ckgate.genpp,v 1.15 2006/06/21 06:18:22 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module PREICGX0P5BA10TR (ECK, E, SE, CK);
output ECK;
input  E, SE, CK;
reg NOTIFIER;

supply1 R, S;

  or       I0 (n1, SE, E);
  udp_tlat I1 (n0, n1, CK, R, S, NOTIFIER);
  and      I2 (ECK, n0, CK);
  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SE$ECK   = 1.0,
      tphl$SE$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SE$CK  = 1.0,
      thold$SE$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      if (E==1'b0 && SE==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b0 && SE==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SE==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SE==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SE == 0), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (SE == 0), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
    $setuphold(posedge CK, posedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER);
    $setuphold(posedge CK, negedge SE, tsetup$SE$CK, thold$SE$CK, NOTIFIER);
  endspecify

endmodule //PREICGX0P5BA10TR
`endcelldefine
//$Id: ckgate.genpp,v 1.15 2006/06/21 06:18:22 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module POSTICGX9BA10TR (ECK, E, SEN, CK);
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, NOTIFIER);
  and      I2 (ECK, n0, CK);
  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SEN$ECK   = 1.0,
      tphl$SEN$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SEN$CK  = 1.0,
      thold$SEN$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      if (E==1'b0 && SEN==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b0 && SEN==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SEN==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SEN==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SEN == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (SEN == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
  endspecify

endmodule //POSTICGX9BA10TR
`endcelldefine
//$Id: ckgate.genpp,v 1.15 2006/06/21 06:18:22 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module POSTICGX7P5BA10TR (ECK, E, SEN, CK);
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, NOTIFIER);
  and      I2 (ECK, n0, CK);
  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SEN$ECK   = 1.0,
      tphl$SEN$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SEN$CK  = 1.0,
      thold$SEN$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      if (E==1'b0 && SEN==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b0 && SEN==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SEN==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SEN==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SEN == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (SEN == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
  endspecify

endmodule //POSTICGX7P5BA10TR
`endcelldefine
//$Id: ckgate.genpp,v 1.15 2006/06/21 06:18:22 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module POSTICGX6BA10TR (ECK, E, SEN, CK);
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, NOTIFIER);
  and      I2 (ECK, n0, CK);
  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SEN$ECK   = 1.0,
      tphl$SEN$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SEN$CK  = 1.0,
      thold$SEN$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      if (E==1'b0 && SEN==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b0 && SEN==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SEN==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SEN==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SEN == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (SEN == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
  endspecify

endmodule //POSTICGX6BA10TR
`endcelldefine
//$Id: ckgate.genpp,v 1.15 2006/06/21 06:18:22 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module POSTICGX5BA10TR (ECK, E, SEN, CK);
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, NOTIFIER);
  and      I2 (ECK, n0, CK);
  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SEN$ECK   = 1.0,
      tphl$SEN$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SEN$CK  = 1.0,
      thold$SEN$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      if (E==1'b0 && SEN==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b0 && SEN==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SEN==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SEN==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SEN == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (SEN == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
  endspecify

endmodule //POSTICGX5BA10TR
`endcelldefine
//$Id: ckgate.genpp,v 1.15 2006/06/21 06:18:22 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module POSTICGX4BA10TR (ECK, E, SEN, CK);
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, NOTIFIER);
  and      I2 (ECK, n0, CK);
  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SEN$ECK   = 1.0,
      tphl$SEN$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SEN$CK  = 1.0,
      thold$SEN$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      if (E==1'b0 && SEN==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b0 && SEN==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SEN==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SEN==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SEN == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (SEN == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
  endspecify

endmodule //POSTICGX4BA10TR
`endcelldefine
//$Id: ckgate.genpp,v 1.15 2006/06/21 06:18:22 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module POSTICGX3P5BA10TR (ECK, E, SEN, CK);
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, NOTIFIER);
  and      I2 (ECK, n0, CK);
  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SEN$ECK   = 1.0,
      tphl$SEN$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SEN$CK  = 1.0,
      thold$SEN$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      if (E==1'b0 && SEN==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b0 && SEN==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SEN==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SEN==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SEN == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (SEN == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
  endspecify

endmodule //POSTICGX3P5BA10TR
`endcelldefine
//$Id: ckgate.genpp,v 1.15 2006/06/21 06:18:22 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module POSTICGX3BA10TR (ECK, E, SEN, CK);
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, NOTIFIER);
  and      I2 (ECK, n0, CK);
  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SEN$ECK   = 1.0,
      tphl$SEN$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SEN$CK  = 1.0,
      thold$SEN$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      if (E==1'b0 && SEN==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b0 && SEN==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SEN==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SEN==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SEN == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (SEN == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
  endspecify

endmodule //POSTICGX3BA10TR
`endcelldefine
//$Id: ckgate.genpp,v 1.15 2006/06/21 06:18:22 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module POSTICGX2P5BA10TR (ECK, E, SEN, CK);
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, NOTIFIER);
  and      I2 (ECK, n0, CK);
  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SEN$ECK   = 1.0,
      tphl$SEN$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SEN$CK  = 1.0,
      thold$SEN$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      if (E==1'b0 && SEN==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b0 && SEN==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SEN==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SEN==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SEN == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (SEN == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
  endspecify

endmodule //POSTICGX2P5BA10TR
`endcelldefine
//$Id: ckgate.genpp,v 1.15 2006/06/21 06:18:22 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module POSTICGX2BA10TR (ECK, E, SEN, CK);
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, NOTIFIER);
  and      I2 (ECK, n0, CK);
  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SEN$ECK   = 1.0,
      tphl$SEN$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SEN$CK  = 1.0,
      thold$SEN$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      if (E==1'b0 && SEN==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b0 && SEN==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SEN==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SEN==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SEN == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (SEN == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
  endspecify

endmodule //POSTICGX2BA10TR
`endcelldefine
//$Id: ckgate.genpp,v 1.15 2006/06/21 06:18:22 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module POSTICGX1P7BA10TR (ECK, E, SEN, CK);
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, NOTIFIER);
  and      I2 (ECK, n0, CK);
  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SEN$ECK   = 1.0,
      tphl$SEN$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SEN$CK  = 1.0,
      thold$SEN$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      if (E==1'b0 && SEN==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b0 && SEN==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SEN==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SEN==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SEN == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (SEN == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
  endspecify

endmodule //POSTICGX1P7BA10TR
`endcelldefine
//$Id: ckgate.genpp,v 1.15 2006/06/21 06:18:22 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module POSTICGX1P4BA10TR (ECK, E, SEN, CK);
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, NOTIFIER);
  and      I2 (ECK, n0, CK);
  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SEN$ECK   = 1.0,
      tphl$SEN$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SEN$CK  = 1.0,
      thold$SEN$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      if (E==1'b0 && SEN==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b0 && SEN==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SEN==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SEN==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SEN == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (SEN == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
  endspecify

endmodule //POSTICGX1P4BA10TR
`endcelldefine
//$Id: ckgate.genpp,v 1.15 2006/06/21 06:18:22 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module POSTICGX1P2BA10TR (ECK, E, SEN, CK);
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, NOTIFIER);
  and      I2 (ECK, n0, CK);
  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SEN$ECK   = 1.0,
      tphl$SEN$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SEN$CK  = 1.0,
      thold$SEN$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      if (E==1'b0 && SEN==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b0 && SEN==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SEN==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SEN==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SEN == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (SEN == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
  endspecify

endmodule //POSTICGX1P2BA10TR
`endcelldefine
//$Id: ckgate.genpp,v 1.15 2006/06/21 06:18:22 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module POSTICGX1BA10TR (ECK, E, SEN, CK);
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, NOTIFIER);
  and      I2 (ECK, n0, CK);
  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SEN$ECK   = 1.0,
      tphl$SEN$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SEN$CK  = 1.0,
      thold$SEN$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      if (E==1'b0 && SEN==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b0 && SEN==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SEN==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SEN==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SEN == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (SEN == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
  endspecify

endmodule //POSTICGX1BA10TR
`endcelldefine
//$Id: ckgate.genpp,v 1.15 2006/06/21 06:18:22 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module POSTICGX16BA10TR (ECK, E, SEN, CK);
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, NOTIFIER);
  and      I2 (ECK, n0, CK);
  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SEN$ECK   = 1.0,
      tphl$SEN$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SEN$CK  = 1.0,
      thold$SEN$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      if (E==1'b0 && SEN==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b0 && SEN==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SEN==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SEN==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SEN == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (SEN == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
  endspecify

endmodule //POSTICGX16BA10TR
`endcelldefine
//$Id: ckgate.genpp,v 1.15 2006/06/21 06:18:22 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module POSTICGX13BA10TR (ECK, E, SEN, CK);
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, NOTIFIER);
  and      I2 (ECK, n0, CK);
  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SEN$ECK   = 1.0,
      tphl$SEN$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SEN$CK  = 1.0,
      thold$SEN$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      if (E==1'b0 && SEN==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b0 && SEN==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SEN==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SEN==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SEN == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (SEN == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
  endspecify

endmodule //POSTICGX13BA10TR
`endcelldefine
//$Id: ckgate.genpp,v 1.15 2006/06/21 06:18:22 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module POSTICGX11BA10TR (ECK, E, SEN, CK);
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, NOTIFIER);
  and      I2 (ECK, n0, CK);
  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SEN$ECK   = 1.0,
      tphl$SEN$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SEN$CK  = 1.0,
      thold$SEN$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      if (E==1'b0 && SEN==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b0 && SEN==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SEN==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SEN==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SEN == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (SEN == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
  endspecify

endmodule //POSTICGX11BA10TR
`endcelldefine
//$Id: ckgate.genpp,v 1.15 2006/06/21 06:18:22 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module POSTICGX0P8BA10TR (ECK, E, SEN, CK);
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, NOTIFIER);
  and      I2 (ECK, n0, CK);
  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SEN$ECK   = 1.0,
      tphl$SEN$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SEN$CK  = 1.0,
      thold$SEN$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      if (E==1'b0 && SEN==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b0 && SEN==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SEN==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SEN==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SEN == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (SEN == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
  endspecify

endmodule //POSTICGX0P8BA10TR
`endcelldefine
//$Id: ckgate.genpp,v 1.15 2006/06/21 06:18:22 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module POSTICGX0P7BA10TR (ECK, E, SEN, CK);
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, NOTIFIER);
  and      I2 (ECK, n0, CK);
  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SEN$ECK   = 1.0,
      tphl$SEN$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SEN$CK  = 1.0,
      thold$SEN$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      if (E==1'b0 && SEN==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b0 && SEN==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SEN==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SEN==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SEN == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (SEN == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
  endspecify

endmodule //POSTICGX0P7BA10TR
`endcelldefine
//$Id: ckgate.genpp,v 1.15 2006/06/21 06:18:22 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module POSTICGX0P6BA10TR (ECK, E, SEN, CK);
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, NOTIFIER);
  and      I2 (ECK, n0, CK);
  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SEN$ECK   = 1.0,
      tphl$SEN$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SEN$CK  = 1.0,
      thold$SEN$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      if (E==1'b0 && SEN==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b0 && SEN==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SEN==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SEN==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SEN == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (SEN == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
  endspecify

endmodule //POSTICGX0P6BA10TR
`endcelldefine
//$Id: ckgate.genpp,v 1.15 2006/06/21 06:18:22 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module POSTICGX0P5BA10TR (ECK, E, SEN, CK);
output ECK;
input  E, SEN, CK;
reg NOTIFIER;

supply1 R, S;

  not      I0 (ovrd, SEN);
  udp_plat I1 (n0, ovrd, CK, E, NOTIFIER);
  and      I2 (ECK, n0, CK);
  specify
    specparam 
      tplh$E$ECK    = 1.0,
      tphl$E$ECK    = 1.0,
      tplh$SEN$ECK   = 1.0,
      tphl$SEN$ECK   = 1.0,
      tplh$CK$ECK   = 1.0,
      tphl$CK$ECK   = 1.0,
      tsetup$E$CK   = 1.0,
      thold$E$CK    = 0.5,
      tsetup$SEN$CK  = 1.0,
      thold$SEN$CK   = 0.5,
      tminpwl$CK    = 1.0,
      tperiod$CK    = 1.0;

    // path delays
      if (E==1'b0 && SEN==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b0 && SEN==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SEN==1'b0) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);
      if (E==1'b1 && SEN==1'b1) (CK *> ECK) = (tplh$CK$ECK,    tphl$CK$ECK);

    // timing checks
    $setuphold(posedge CK &&& (SEN == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (SEN == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $width(negedge CK, tminpwl$CK, 0, NOTIFIER);
    $period(negedge CK, tperiod$CK, NOTIFIER);
  endspecify

endmodule //POSTICGX0P5BA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR6X6MA10TR (Y, A, B, C, D, E, F);
output Y;
input A, B, C, D, E, F;

  or (Y, A, B, C, D, E, F);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0,
      tplh$E$Y = 1.0,
      tphl$E$Y = 1.0,
      tplh$F$Y = 1.0,
      tphl$F$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
    (E *> Y) = (tplh$E$Y, tphl$E$Y);
    (F *> Y) = (tplh$F$Y, tphl$F$Y);
  endspecify
endmodule // OR6X6MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR6X4MA10TR (Y, A, B, C, D, E, F);
output Y;
input A, B, C, D, E, F;

  or (Y, A, B, C, D, E, F);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0,
      tplh$E$Y = 1.0,
      tphl$E$Y = 1.0,
      tplh$F$Y = 1.0,
      tphl$F$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
    (E *> Y) = (tplh$E$Y, tphl$E$Y);
    (F *> Y) = (tplh$F$Y, tphl$F$Y);
  endspecify
endmodule // OR6X4MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR6X3MA10TR (Y, A, B, C, D, E, F);
output Y;
input A, B, C, D, E, F;

  or (Y, A, B, C, D, E, F);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0,
      tplh$E$Y = 1.0,
      tphl$E$Y = 1.0,
      tplh$F$Y = 1.0,
      tphl$F$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
    (E *> Y) = (tplh$E$Y, tphl$E$Y);
    (F *> Y) = (tplh$F$Y, tphl$F$Y);
  endspecify
endmodule // OR6X3MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR6X2MA10TR (Y, A, B, C, D, E, F);
output Y;
input A, B, C, D, E, F;

  or (Y, A, B, C, D, E, F);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0,
      tplh$E$Y = 1.0,
      tphl$E$Y = 1.0,
      tplh$F$Y = 1.0,
      tphl$F$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
    (E *> Y) = (tplh$E$Y, tphl$E$Y);
    (F *> Y) = (tplh$F$Y, tphl$F$Y);
  endspecify
endmodule // OR6X2MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR6X1P4MA10TR (Y, A, B, C, D, E, F);
output Y;
input A, B, C, D, E, F;

  or (Y, A, B, C, D, E, F);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0,
      tplh$E$Y = 1.0,
      tphl$E$Y = 1.0,
      tplh$F$Y = 1.0,
      tphl$F$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
    (E *> Y) = (tplh$E$Y, tphl$E$Y);
    (F *> Y) = (tplh$F$Y, tphl$F$Y);
  endspecify
endmodule // OR6X1P4MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR6X1MA10TR (Y, A, B, C, D, E, F);
output Y;
input A, B, C, D, E, F;

  or (Y, A, B, C, D, E, F);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0,
      tplh$E$Y = 1.0,
      tphl$E$Y = 1.0,
      tplh$F$Y = 1.0,
      tphl$F$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
    (E *> Y) = (tplh$E$Y, tphl$E$Y);
    (F *> Y) = (tplh$F$Y, tphl$F$Y);
  endspecify
endmodule // OR6X1MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR6X0P7MA10TR (Y, A, B, C, D, E, F);
output Y;
input A, B, C, D, E, F;

  or (Y, A, B, C, D, E, F);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0,
      tplh$E$Y = 1.0,
      tphl$E$Y = 1.0,
      tplh$F$Y = 1.0,
      tphl$F$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
    (E *> Y) = (tplh$E$Y, tphl$E$Y);
    (F *> Y) = (tplh$F$Y, tphl$F$Y);
  endspecify
endmodule // OR6X0P7MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR6X0P5MA10TR (Y, A, B, C, D, E, F);
output Y;
input A, B, C, D, E, F;

  or (Y, A, B, C, D, E, F);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0,
      tplh$E$Y = 1.0,
      tphl$E$Y = 1.0,
      tplh$F$Y = 1.0,
      tphl$F$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
    (E *> Y) = (tplh$E$Y, tphl$E$Y);
    (F *> Y) = (tplh$F$Y, tphl$F$Y);
  endspecify
endmodule // OR6X0P5MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR4X8MA10TR (Y, A, B, C, D);
output Y;
input A, B, C, D;

  or (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // OR4X8MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR4X6MA10TR (Y, A, B, C, D);
output Y;
input A, B, C, D;

  or (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // OR4X6MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR4X4MA10TR (Y, A, B, C, D);
output Y;
input A, B, C, D;

  or (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // OR4X4MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR4X3MA10TR (Y, A, B, C, D);
output Y;
input A, B, C, D;

  or (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // OR4X3MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR4X2MA10TR (Y, A, B, C, D);
output Y;
input A, B, C, D;

  or (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // OR4X2MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR4X1P4MA10TR (Y, A, B, C, D);
output Y;
input A, B, C, D;

  or (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // OR4X1P4MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR4X1MA10TR (Y, A, B, C, D);
output Y;
input A, B, C, D;

  or (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // OR4X1MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR4X0P7MA10TR (Y, A, B, C, D);
output Y;
input A, B, C, D;

  or (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // OR4X0P7MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR4X0P5MA10TR (Y, A, B, C, D);
output Y;
input A, B, C, D;

  or (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // OR4X0P5MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR3X8MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  or (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // OR3X8MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR3X6MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  or (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // OR3X6MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR3X4MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  or (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // OR3X4MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR3X3MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  or (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // OR3X3MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR3X2MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  or (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // OR3X2MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR3X1P4MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  or (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // OR3X1P4MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR3X1MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  or (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // OR3X1MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR3X0P7MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  or (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // OR3X0P7MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR3X0P5MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  or (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // OR3X0P5MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR2X8MA10TR (Y, A, B);
output Y;
input A, B;

  or (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // OR2X8MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR2X6MA10TR (Y, A, B);
output Y;
input A, B;

  or (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // OR2X6MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR2X4MA10TR (Y, A, B);
output Y;
input A, B;

  or (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // OR2X4MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR2X3MA10TR (Y, A, B);
output Y;
input A, B;

  or (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // OR2X3MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR2X2MA10TR (Y, A, B);
output Y;
input A, B;

  or (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // OR2X2MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR2X1P4MA10TR (Y, A, B);
output Y;
input A, B;

  or (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // OR2X1P4MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR2X1MA10TR (Y, A, B);
output Y;
input A, B;

  or (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // OR2X1MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR2X11MA10TR (Y, A, B);
output Y;
input A, B;

  or (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // OR2X11MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR2X0P7MA10TR (Y, A, B);
output Y;
input A, B;

  or (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // OR2X0P7MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OR2X0P5MA10TR (Y, A, B);
output Y;
input A, B;

  or (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // OR2X0P5MA10TR
`endcelldefine
//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI2XB1X8MA10TR (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;

  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);
    if (A0 == 1'b0 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OAI2XB1X8MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI2XB1X6MA10TR (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;

  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);
    if (A0 == 1'b0 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OAI2XB1X6MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI2XB1X4MA10TR (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;

  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);
    if (A0 == 1'b0 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OAI2XB1X4MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI2XB1X3MA10TR (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;

  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);
    if (A0 == 1'b0 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OAI2XB1X3MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI2XB1X2MA10TR (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;

  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);
    if (A0 == 1'b0 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OAI2XB1X2MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI2XB1X1P4MA10TR (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;

  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);
    if (A0 == 1'b0 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OAI2XB1X1P4MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI2XB1X1MA10TR (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;

  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);
    if (A0 == 1'b0 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OAI2XB1X1MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI2XB1X0P7MA10TR (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;

  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);
    if (A0 == 1'b0 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OAI2XB1X0P7MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI2XB1X0P5MA10TR (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;

  not  I0 (outA1, A1N);
  or   I1 (outA, A0, outA1);
  nand I2 (Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);
    if (A0 == 1'b0 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OAI2XB1X0P5MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI22X8MA10TR (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // OAI22X8MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI22X6MA10TR (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // OAI22X6MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI22X4MA10TR (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // OAI22X4MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI22X3MA10TR (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // OAI22X3MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI22X2MA10TR (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // OAI22X2MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI22X1P4MA10TR (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // OAI22X1P4MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI22X1MA10TR (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // OAI22X1MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI22X0P7MA10TR (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // OAI22X0P7MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI22X0P5MA10TR (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // OAI22X0P5MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI222X4MA10TR (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand I3(Y, outA, outB, outC);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0,
      tplh$C1$Y = 1.0,
      tphl$C1$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y);

  endspecify
endmodule // OAI222X4MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI222X3MA10TR (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand I3(Y, outA, outB, outC);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0,
      tplh$C1$Y = 1.0,
      tphl$C1$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y);

  endspecify
endmodule // OAI222X3MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI222X2MA10TR (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand I3(Y, outA, outB, outC);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0,
      tplh$C1$Y = 1.0,
      tphl$C1$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y);

  endspecify
endmodule // OAI222X2MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI222X1P4MA10TR (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand I3(Y, outA, outB, outC);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0,
      tplh$C1$Y = 1.0,
      tphl$C1$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y);

  endspecify
endmodule // OAI222X1P4MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI222X1MA10TR (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand I3(Y, outA, outB, outC);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0,
      tplh$C1$Y = 1.0,
      tphl$C1$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y);

  endspecify
endmodule // OAI222X1MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI222X0P7MA10TR (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand I3(Y, outA, outB, outC);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0,
      tplh$C1$Y = 1.0,
      tphl$C1$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y);

  endspecify
endmodule // OAI222X0P7MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI222X0P5MA10TR (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  or   I2(outC, C0, C1);
  nand I3(Y, outA, outB, outC);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0,
      tplh$C1$Y = 1.0,
      tphl$C1$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && C1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y);

  endspecify
endmodule // OAI222X0P5MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI221X4MA10TR (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, C0, outB, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && C0 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // OAI221X4MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI221X3MA10TR (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, C0, outB, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && C0 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // OAI221X3MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI221X2MA10TR (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, C0, outB, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && C0 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // OAI221X2MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI221X1P4MA10TR (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, C0, outB, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && C0 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // OAI221X1P4MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI221X1MA10TR (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, C0, outB, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && C0 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // OAI221X1MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI221X0P7MA10TR (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, C0, outB, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && C0 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // OAI221X0P7MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI221X0P5MA10TR (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  nand I2(Y, C0, outB, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && C0 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && C0 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // OAI221X0P5MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI21BX8MA10TR (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;

  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand I2 (Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0N$Y = 1.0,
      tphl$B0N$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0N == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0N == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y);

  endspecify
endmodule // OAI21BX8MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI21BX6MA10TR (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;

  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand I2 (Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0N$Y = 1.0,
      tphl$B0N$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0N == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0N == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y);

  endspecify
endmodule // OAI21BX6MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI21BX4MA10TR (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;

  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand I2 (Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0N$Y = 1.0,
      tphl$B0N$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0N == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0N == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y);

  endspecify
endmodule // OAI21BX4MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI21BX3MA10TR (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;

  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand I2 (Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0N$Y = 1.0,
      tphl$B0N$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0N == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0N == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y);

  endspecify
endmodule // OAI21BX3MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI21BX2MA10TR (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;

  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand I2 (Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0N$Y = 1.0,
      tphl$B0N$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0N == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0N == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y);

  endspecify
endmodule // OAI21BX2MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI21BX1P4MA10TR (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;

  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand I2 (Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0N$Y = 1.0,
      tphl$B0N$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0N == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0N == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y);

  endspecify
endmodule // OAI21BX1P4MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI21BX1MA10TR (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;

  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand I2 (Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0N$Y = 1.0,
      tphl$B0N$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0N == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0N == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y);

  endspecify
endmodule // OAI21BX1MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI21BX0P7MA10TR (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;

  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand I2 (Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0N$Y = 1.0,
      tphl$B0N$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0N == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0N == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y);

  endspecify
endmodule // OAI21BX0P7MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI21BX0P5MA10TR (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;

  not  I0 (outB, B0N);
  or   I1 (outA, A0,  A1);
  nand I2 (Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0N$Y = 1.0,
      tphl$B0N$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0N == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0N == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y);

  endspecify
endmodule // OAI21BX0P5MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI21X8MA10TR (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  or   I0(outA, A0, A1);
  nand I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OAI21X8MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI21X6MA10TR (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  or   I0(outA, A0, A1);
  nand I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OAI21X6MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI21X4MA10TR (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  or   I0(outA, A0, A1);
  nand I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OAI21X4MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI21X3MA10TR (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  or   I0(outA, A0, A1);
  nand I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OAI21X3MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI21X2MA10TR (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  or   I0(outA, A0, A1);
  nand I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OAI21X2MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI21X1P4MA10TR (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  or   I0(outA, A0, A1);
  nand I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OAI21X1P4MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI21X1MA10TR (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  or   I0(outA, A0, A1);
  nand I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OAI21X1MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI21X0P7MA10TR (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  or   I0(outA, A0, A1);
  nand I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OAI21X0P7MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI21X0P5MA10TR (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  or   I0(outA, A0, A1);
  nand I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OAI21X0P5MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI211X4MA10TR (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;

  or   I0(outA, A0, A1);
  nand I1(Y, B0, C0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b0 && A1 == 1'b1 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // OAI211X4MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI211X3MA10TR (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;

  or   I0(outA, A0, A1);
  nand I1(Y, B0, C0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b0 && A1 == 1'b1 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // OAI211X3MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI211X2MA10TR (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;

  or   I0(outA, A0, A1);
  nand I1(Y, B0, C0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b0 && A1 == 1'b1 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // OAI211X2MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI211X1P4MA10TR (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;

  or   I0(outA, A0, A1);
  nand I1(Y, B0, C0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b0 && A1 == 1'b1 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // OAI211X1P4MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI211X1MA10TR (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;

  or   I0(outA, A0, A1);
  nand I1(Y, B0, C0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b0 && A1 == 1'b1 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // OAI211X1MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI211X0P7MA10TR (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;

  or   I0(outA, A0, A1);
  nand I1(Y, B0, C0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b0 && A1 == 1'b1 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // OAI211X0P7MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OAI211X0P5MA10TR (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;

  or   I0(outA, A0, A1);
  nand I1(Y, B0, C0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b0 && A1 == 1'b1 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && C0 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && B0 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // OAI211X0P5MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OA22X8MA10TR (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // OA22X8MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OA22X6MA10TR (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // OA22X6MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OA22X4MA10TR (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // OA22X4MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OA22X3MA10TR (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // OA22X3MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OA22X2MA10TR (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // OA22X2MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OA22X1P4MA10TR (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // OA22X1P4MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OA22X1MA10TR (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // OA22X1MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OA22X0P7MA10TR (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // OA22X0P7MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OA22X0P5MA10TR (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  or   I0(outA, A0, A1);
  or   I1(outB, B0, B1);
  and I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && B0 == 1'b1 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b1 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b0 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // OA22X0P5MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OA21X8MA10TR (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  or   I0(outA, A0, A1);
  and I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OA21X8MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OA21X6MA10TR (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  or   I0(outA, A0, A1);
  and I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OA21X6MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OA21X4MA10TR (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  or   I0(outA, A0, A1);
  and I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OA21X4MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OA21X3MA10TR (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  or   I0(outA, A0, A1);
  and I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OA21X3MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OA21X2MA10TR (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  or   I0(outA, A0, A1);
  and I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OA21X2MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OA21X1P4MA10TR (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  or   I0(outA, A0, A1);
  and I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OA21X1P4MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OA21X1MA10TR (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  or   I0(outA, A0, A1);
  and I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OA21X1MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OA21X0P7MA10TR (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  or   I0(outA, A0, A1);
  and I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OA21X0P7MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OA21X0P5MA10TR (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  or   I0(outA, A0, A1);
  and I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // OA21X0P5MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OA211X6MA10TR (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;

  or   I0(outA, A0, A1);
  and I1(Y, B0, C0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
   if ( A0 == 0 && A1 == 1 && C0 == 1  )
      ( B0 *> Y) = ( tplh$B0$Y, tphl$B0$Y);
   if ( A0 == 1 && A1 == 1 && C0 == 1  )
      ( B0 *> Y) = ( tplh$B0$Y, tphl$B0$Y);
   if ( A0 == 1 && A1 == 0 && C0 == 1  )
      ( B0 *> Y) = ( tplh$B0$Y, tphl$B0$Y);
   if ( A0 == 0 && A1 == 1 && B0 == 1  )
      ( C0 *> Y) = ( tplh$C0$Y, tphl$C0$Y);
   if ( A0 == 1 && A1 == 0 && B0 == 1  )
      ( C0 *> Y) = ( tplh$C0$Y, tphl$C0$Y);
   if ( A0 == 1 && A1 == 1 && B0 == 1  )
      ( C0 *> Y) = ( tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // OA211X6MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OA211X4MA10TR (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;

  or   I0(outA, A0, A1);
  and I1(Y, B0, C0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
   if ( A0 == 0 && A1 == 1 && C0 == 1  )
      ( B0 *> Y) = ( tplh$B0$Y, tphl$B0$Y);
   if ( A0 == 1 && A1 == 1 && C0 == 1  )
      ( B0 *> Y) = ( tplh$B0$Y, tphl$B0$Y);
   if ( A0 == 1 && A1 == 0 && C0 == 1  )
      ( B0 *> Y) = ( tplh$B0$Y, tphl$B0$Y);
   if ( A0 == 0 && A1 == 1 && B0 == 1  )
      ( C0 *> Y) = ( tplh$C0$Y, tphl$C0$Y);
   if ( A0 == 1 && A1 == 0 && B0 == 1  )
      ( C0 *> Y) = ( tplh$C0$Y, tphl$C0$Y);
   if ( A0 == 1 && A1 == 1 && B0 == 1  )
      ( C0 *> Y) = ( tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // OA211X4MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OA211X3MA10TR (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;

  or   I0(outA, A0, A1);
  and I1(Y, B0, C0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
   if ( A0 == 0 && A1 == 1 && C0 == 1  )
      ( B0 *> Y) = ( tplh$B0$Y, tphl$B0$Y);
   if ( A0 == 1 && A1 == 1 && C0 == 1  )
      ( B0 *> Y) = ( tplh$B0$Y, tphl$B0$Y);
   if ( A0 == 1 && A1 == 0 && C0 == 1  )
      ( B0 *> Y) = ( tplh$B0$Y, tphl$B0$Y);
   if ( A0 == 0 && A1 == 1 && B0 == 1  )
      ( C0 *> Y) = ( tplh$C0$Y, tphl$C0$Y);
   if ( A0 == 1 && A1 == 0 && B0 == 1  )
      ( C0 *> Y) = ( tplh$C0$Y, tphl$C0$Y);
   if ( A0 == 1 && A1 == 1 && B0 == 1  )
      ( C0 *> Y) = ( tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // OA211X3MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OA211X2MA10TR (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;

  or   I0(outA, A0, A1);
  and I1(Y, B0, C0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
   if ( A0 == 0 && A1 == 1 && C0 == 1  )
      ( B0 *> Y) = ( tplh$B0$Y, tphl$B0$Y);
   if ( A0 == 1 && A1 == 1 && C0 == 1  )
      ( B0 *> Y) = ( tplh$B0$Y, tphl$B0$Y);
   if ( A0 == 1 && A1 == 0 && C0 == 1  )
      ( B0 *> Y) = ( tplh$B0$Y, tphl$B0$Y);
   if ( A0 == 0 && A1 == 1 && B0 == 1  )
      ( C0 *> Y) = ( tplh$C0$Y, tphl$C0$Y);
   if ( A0 == 1 && A1 == 0 && B0 == 1  )
      ( C0 *> Y) = ( tplh$C0$Y, tphl$C0$Y);
   if ( A0 == 1 && A1 == 1 && B0 == 1  )
      ( C0 *> Y) = ( tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // OA211X2MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OA211X1P4MA10TR (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;

  or   I0(outA, A0, A1);
  and I1(Y, B0, C0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
   if ( A0 == 0 && A1 == 1 && C0 == 1  )
      ( B0 *> Y) = ( tplh$B0$Y, tphl$B0$Y);
   if ( A0 == 1 && A1 == 1 && C0 == 1  )
      ( B0 *> Y) = ( tplh$B0$Y, tphl$B0$Y);
   if ( A0 == 1 && A1 == 0 && C0 == 1  )
      ( B0 *> Y) = ( tplh$B0$Y, tphl$B0$Y);
   if ( A0 == 0 && A1 == 1 && B0 == 1  )
      ( C0 *> Y) = ( tplh$C0$Y, tphl$C0$Y);
   if ( A0 == 1 && A1 == 0 && B0 == 1  )
      ( C0 *> Y) = ( tplh$C0$Y, tphl$C0$Y);
   if ( A0 == 1 && A1 == 1 && B0 == 1  )
      ( C0 *> Y) = ( tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // OA211X1P4MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OA211X1MA10TR (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;

  or   I0(outA, A0, A1);
  and I1(Y, B0, C0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
   if ( A0 == 0 && A1 == 1 && C0 == 1  )
      ( B0 *> Y) = ( tplh$B0$Y, tphl$B0$Y);
   if ( A0 == 1 && A1 == 1 && C0 == 1  )
      ( B0 *> Y) = ( tplh$B0$Y, tphl$B0$Y);
   if ( A0 == 1 && A1 == 0 && C0 == 1  )
      ( B0 *> Y) = ( tplh$B0$Y, tphl$B0$Y);
   if ( A0 == 0 && A1 == 1 && B0 == 1  )
      ( C0 *> Y) = ( tplh$C0$Y, tphl$C0$Y);
   if ( A0 == 1 && A1 == 0 && B0 == 1  )
      ( C0 *> Y) = ( tplh$C0$Y, tphl$C0$Y);
   if ( A0 == 1 && A1 == 1 && B0 == 1  )
      ( C0 *> Y) = ( tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // OA211X1MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OA211X0P7MA10TR (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;

  or   I0(outA, A0, A1);
  and I1(Y, B0, C0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
   if ( A0 == 0 && A1 == 1 && C0 == 1  )
      ( B0 *> Y) = ( tplh$B0$Y, tphl$B0$Y);
   if ( A0 == 1 && A1 == 1 && C0 == 1  )
      ( B0 *> Y) = ( tplh$B0$Y, tphl$B0$Y);
   if ( A0 == 1 && A1 == 0 && C0 == 1  )
      ( B0 *> Y) = ( tplh$B0$Y, tphl$B0$Y);
   if ( A0 == 0 && A1 == 1 && B0 == 1  )
      ( C0 *> Y) = ( tplh$C0$Y, tphl$C0$Y);
   if ( A0 == 1 && A1 == 0 && B0 == 1  )
      ( C0 *> Y) = ( tplh$C0$Y, tphl$C0$Y);
   if ( A0 == 1 && A1 == 1 && B0 == 1  )
      ( C0 *> Y) = ( tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // OA211X0P7MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module OA211X0P5MA10TR (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;

  or   I0(outA, A0, A1);
  and I1(Y, B0, C0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
   if ( A0 == 0 && A1 == 1 && C0 == 1  )
      ( B0 *> Y) = ( tplh$B0$Y, tphl$B0$Y);
   if ( A0 == 1 && A1 == 1 && C0 == 1  )
      ( B0 *> Y) = ( tplh$B0$Y, tphl$B0$Y);
   if ( A0 == 1 && A1 == 0 && C0 == 1  )
      ( B0 *> Y) = ( tplh$B0$Y, tphl$B0$Y);
   if ( A0 == 0 && A1 == 1 && B0 == 1  )
      ( C0 *> Y) = ( tplh$C0$Y, tphl$C0$Y);
   if ( A0 == 1 && A1 == 0 && B0 == 1  )
      ( C0 *> Y) = ( tplh$C0$Y, tphl$C0$Y);
   if ( A0 == 1 && A1 == 1 && B0 == 1  )
      ( C0 *> Y) = ( tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // OA211X0P5MA10TR
`endcelldefine





//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR3X4MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  nor (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NOR3X4MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR3X4AA10TR (Y, A, B, C);
output Y;
input A, B, C;

  nor (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NOR3X4AA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR3X3MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  nor (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NOR3X3MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR3X3AA10TR (Y, A, B, C);
output Y;
input A, B, C;

  nor (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NOR3X3AA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR3X2MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  nor (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NOR3X2MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR3X2AA10TR (Y, A, B, C);
output Y;
input A, B, C;

  nor (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NOR3X2AA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR3X1P4MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  nor (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NOR3X1P4MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR3X1P4AA10TR (Y, A, B, C);
output Y;
input A, B, C;

  nor (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NOR3X1P4AA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR3X1MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  nor (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NOR3X1MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR3X1AA10TR (Y, A, B, C);
output Y;
input A, B, C;

  nor (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NOR3X1AA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR3X0P7MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  nor (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NOR3X0P7MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR3X0P7AA10TR (Y, A, B, C);
output Y;
input A, B, C;

  nor (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NOR3X0P7AA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR3X0P5MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  nor (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NOR3X0P5MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR3X0P5AA10TR (Y, A, B, C);
output Y;
input A, B, C;

  nor (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NOR3X0P5AA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2XBX8MA10TR (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nor (Y, A, Bx);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$BN$Y = 1.0,
      tphl$BN$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (BN *> Y) = (tplh$BN$Y, tphl$BN$Y);
  endspecify
endmodule // NOR2XBX8MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2XBX6MA10TR (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nor (Y, A, Bx);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$BN$Y = 1.0,
      tphl$BN$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (BN *> Y) = (tplh$BN$Y, tphl$BN$Y);
  endspecify
endmodule // NOR2XBX6MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2XBX4MA10TR (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nor (Y, A, Bx);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$BN$Y = 1.0,
      tphl$BN$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (BN *> Y) = (tplh$BN$Y, tphl$BN$Y);
  endspecify
endmodule // NOR2XBX4MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2XBX3MA10TR (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nor (Y, A, Bx);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$BN$Y = 1.0,
      tphl$BN$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (BN *> Y) = (tplh$BN$Y, tphl$BN$Y);
  endspecify
endmodule // NOR2XBX3MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2XBX2MA10TR (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nor (Y, A, Bx);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$BN$Y = 1.0,
      tphl$BN$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (BN *> Y) = (tplh$BN$Y, tphl$BN$Y);
  endspecify
endmodule // NOR2XBX2MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2XBX1P4MA10TR (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nor (Y, A, Bx);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$BN$Y = 1.0,
      tphl$BN$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (BN *> Y) = (tplh$BN$Y, tphl$BN$Y);
  endspecify
endmodule // NOR2XBX1P4MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2XBX1MA10TR (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nor (Y, A, Bx);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$BN$Y = 1.0,
      tphl$BN$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (BN *> Y) = (tplh$BN$Y, tphl$BN$Y);
  endspecify
endmodule // NOR2XBX1MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2XBX0P7MA10TR (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nor (Y, A, Bx);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$BN$Y = 1.0,
      tphl$BN$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (BN *> Y) = (tplh$BN$Y, tphl$BN$Y);
  endspecify
endmodule // NOR2XBX0P7MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2XBX0P5MA10TR (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nor (Y, A, Bx);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$BN$Y = 1.0,
      tphl$BN$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (BN *> Y) = (tplh$BN$Y, tphl$BN$Y);
  endspecify
endmodule // NOR2XBX0P5MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2BX8MA10TR (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nor (Y, Ax, B);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NOR2BX8MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2BX6MA10TR (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nor (Y, Ax, B);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NOR2BX6MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2BX4MA10TR (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nor (Y, Ax, B);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NOR2BX4MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2BX3MA10TR (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nor (Y, Ax, B);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NOR2BX3MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2BX2MA10TR (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nor (Y, Ax, B);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NOR2BX2MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2BX1P4MA10TR (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nor (Y, Ax, B);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NOR2BX1P4MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2BX1MA10TR (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nor (Y, Ax, B);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NOR2BX1MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2BX0P7MA10TR (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nor (Y, Ax, B);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NOR2BX0P7MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2BX0P5MA10TR (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nor (Y, Ax, B);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NOR2BX0P5MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2X8MA10TR (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NOR2X8MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2X8AA10TR (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NOR2X8AA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2X6MA10TR (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NOR2X6MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2X6AA10TR (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NOR2X6AA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2X4MA10TR (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NOR2X4MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2X4AA10TR (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NOR2X4AA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2X3MA10TR (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NOR2X3MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2X3AA10TR (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NOR2X3AA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2X2MA10TR (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NOR2X2MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2X2AA10TR (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NOR2X2AA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2X1P4MA10TR (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NOR2X1P4MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2X1P4AA10TR (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NOR2X1P4AA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2X1MA10TR (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NOR2X1MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2X1AA10TR (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NOR2X1AA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2X0P7MA10TR (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NOR2X0P7MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2X0P7AA10TR (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NOR2X0P7AA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2X0P5MA10TR (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NOR2X0P5MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NOR2X0P5AA10TR (Y, A, B);
output Y;
input A, B;

  nor (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NOR2X0P5AA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND4XXXBX4MA10TR (Y, A, B, C, DN);
output Y;
input A, B, C, DN;

  not (Dx, DN);
  nand (Y, A, B, C, Dx);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$DN$Y = 1.0,
      tphl$DN$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (DN *> Y) = (tplh$DN$Y, tphl$DN$Y);
  endspecify
endmodule // NAND4XXXBX4MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND4XXXBX3MA10TR (Y, A, B, C, DN);
output Y;
input A, B, C, DN;

  not (Dx, DN);
  nand (Y, A, B, C, Dx);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$DN$Y = 1.0,
      tphl$DN$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (DN *> Y) = (tplh$DN$Y, tphl$DN$Y);
  endspecify
endmodule // NAND4XXXBX3MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND4XXXBX2MA10TR (Y, A, B, C, DN);
output Y;
input A, B, C, DN;

  not (Dx, DN);
  nand (Y, A, B, C, Dx);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$DN$Y = 1.0,
      tphl$DN$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (DN *> Y) = (tplh$DN$Y, tphl$DN$Y);
  endspecify
endmodule // NAND4XXXBX2MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND4XXXBX1P4MA10TR (Y, A, B, C, DN);
output Y;
input A, B, C, DN;

  not (Dx, DN);
  nand (Y, A, B, C, Dx);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$DN$Y = 1.0,
      tphl$DN$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (DN *> Y) = (tplh$DN$Y, tphl$DN$Y);
  endspecify
endmodule // NAND4XXXBX1P4MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND4XXXBX1MA10TR (Y, A, B, C, DN);
output Y;
input A, B, C, DN;

  not (Dx, DN);
  nand (Y, A, B, C, Dx);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$DN$Y = 1.0,
      tphl$DN$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (DN *> Y) = (tplh$DN$Y, tphl$DN$Y);
  endspecify
endmodule // NAND4XXXBX1MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND4XXXBX0P7MA10TR (Y, A, B, C, DN);
output Y;
input A, B, C, DN;

  not (Dx, DN);
  nand (Y, A, B, C, Dx);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$DN$Y = 1.0,
      tphl$DN$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (DN *> Y) = (tplh$DN$Y, tphl$DN$Y);
  endspecify
endmodule // NAND4XXXBX0P7MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND4XXXBX0P5MA10TR (Y, A, B, C, DN);
output Y;
input A, B, C, DN;

  not (Dx, DN);
  nand (Y, A, B, C, Dx);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$DN$Y = 1.0,
      tphl$DN$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (DN *> Y) = (tplh$DN$Y, tphl$DN$Y);
  endspecify
endmodule // NAND4XXXBX0P5MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND4BX4MA10TR (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand (Y, Ax, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NAND4BX4MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND4BX3MA10TR (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand (Y, Ax, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NAND4BX3MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND4BX2MA10TR (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand (Y, Ax, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NAND4BX2MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND4BX1P4MA10TR (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand (Y, Ax, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NAND4BX1P4MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND4BX1MA10TR (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand (Y, Ax, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NAND4BX1MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND4BX0P7MA10TR (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand (Y, Ax, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NAND4BX0P7MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND4BX0P5MA10TR (Y, AN, B, C, D);
output Y;
input AN, B, C, D;

  not (Ax, AN);
  nand (Y, Ax, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NAND4BX0P5MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND4X4MA10TR (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NAND4X4MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND4X4AA10TR (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NAND4X4AA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND4X3MA10TR (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NAND4X3MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND4X3AA10TR (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NAND4X3AA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND4X2MA10TR (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NAND4X2MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND4X2AA10TR (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NAND4X2AA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND4X1P4MA10TR (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NAND4X1P4MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND4X1P4AA10TR (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NAND4X1P4AA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND4X1MA10TR (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NAND4X1MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND4X1AA10TR (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NAND4X1AA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND4X0P7MA10TR (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NAND4X0P7MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND4X0P7AA10TR (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NAND4X0P7AA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND4X0P5MA10TR (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NAND4X0P5MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND4X0P5AA10TR (Y, A, B, C, D);
output Y;
input A, B, C, D;

  nand (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // NAND4X0P5AA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND3XXBX6MA10TR (Y, A, B, CN);
output Y;
input A, B, CN;

  not (Cx, CN);
  nand (Y, A, B, Cx);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$CN$Y = 1.0,
      tphl$CN$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (CN *> Y) = (tplh$CN$Y, tphl$CN$Y);
  endspecify
endmodule // NAND3XXBX6MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND3XXBX4MA10TR (Y, A, B, CN);
output Y;
input A, B, CN;

  not (Cx, CN);
  nand (Y, A, B, Cx);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$CN$Y = 1.0,
      tphl$CN$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (CN *> Y) = (tplh$CN$Y, tphl$CN$Y);
  endspecify
endmodule // NAND3XXBX4MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND3XXBX3MA10TR (Y, A, B, CN);
output Y;
input A, B, CN;

  not (Cx, CN);
  nand (Y, A, B, Cx);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$CN$Y = 1.0,
      tphl$CN$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (CN *> Y) = (tplh$CN$Y, tphl$CN$Y);
  endspecify
endmodule // NAND3XXBX3MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND3XXBX2MA10TR (Y, A, B, CN);
output Y;
input A, B, CN;

  not (Cx, CN);
  nand (Y, A, B, Cx);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$CN$Y = 1.0,
      tphl$CN$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (CN *> Y) = (tplh$CN$Y, tphl$CN$Y);
  endspecify
endmodule // NAND3XXBX2MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND3XXBX1P4MA10TR (Y, A, B, CN);
output Y;
input A, B, CN;

  not (Cx, CN);
  nand (Y, A, B, Cx);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$CN$Y = 1.0,
      tphl$CN$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (CN *> Y) = (tplh$CN$Y, tphl$CN$Y);
  endspecify
endmodule // NAND3XXBX1P4MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND3XXBX1MA10TR (Y, A, B, CN);
output Y;
input A, B, CN;

  not (Cx, CN);
  nand (Y, A, B, Cx);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$CN$Y = 1.0,
      tphl$CN$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (CN *> Y) = (tplh$CN$Y, tphl$CN$Y);
  endspecify
endmodule // NAND3XXBX1MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND3XXBX0P7MA10TR (Y, A, B, CN);
output Y;
input A, B, CN;

  not (Cx, CN);
  nand (Y, A, B, Cx);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$CN$Y = 1.0,
      tphl$CN$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (CN *> Y) = (tplh$CN$Y, tphl$CN$Y);
  endspecify
endmodule // NAND3XXBX0P7MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND3XXBX0P5MA10TR (Y, A, B, CN);
output Y;
input A, B, CN;

  not (Cx, CN);
  nand (Y, A, B, Cx);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$CN$Y = 1.0,
      tphl$CN$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (CN *> Y) = (tplh$CN$Y, tphl$CN$Y);
  endspecify
endmodule // NAND3XXBX0P5MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND3BX6MA10TR (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nand (Y, Ax, B, C);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NAND3BX6MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND3BX4MA10TR (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nand (Y, Ax, B, C);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NAND3BX4MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND3BX3MA10TR (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nand (Y, Ax, B, C);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NAND3BX3MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND3BX2MA10TR (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nand (Y, Ax, B, C);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NAND3BX2MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND3BX1P4MA10TR (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nand (Y, Ax, B, C);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NAND3BX1P4MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND3BX1MA10TR (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nand (Y, Ax, B, C);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NAND3BX1MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND3BX0P7MA10TR (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nand (Y, Ax, B, C);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NAND3BX0P7MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND3BX0P5MA10TR (Y, AN, B, C);
output Y;
input AN, B, C;

  not (Ax, AN);
  nand (Y, Ax, B, C);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NAND3BX0P5MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND3X6MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NAND3X6MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND3X6AA10TR (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NAND3X6AA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND3X4MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NAND3X4MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND3X4AA10TR (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NAND3X4AA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND3X3MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NAND3X3MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND3X3AA10TR (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NAND3X3AA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND3X2MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NAND3X2MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND3X2AA10TR (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NAND3X2AA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND3X1P4MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NAND3X1P4MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND3X1P4AA10TR (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NAND3X1P4AA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND3X1MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NAND3X1MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND3X1AA10TR (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NAND3X1AA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND3X0P7MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NAND3X0P7MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND3X0P7AA10TR (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NAND3X0P7AA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND3X0P5MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NAND3X0P5MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND3X0P5AA10TR (Y, A, B, C);
output Y;
input A, B, C;

  nand (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // NAND3X0P5AA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2XBX8MA10TR (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nand (Y, A, Bx);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$BN$Y = 1.0,
      tphl$BN$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (BN *> Y) = (tplh$BN$Y, tphl$BN$Y);
  endspecify
endmodule // NAND2XBX8MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2XBX6MA10TR (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nand (Y, A, Bx);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$BN$Y = 1.0,
      tphl$BN$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (BN *> Y) = (tplh$BN$Y, tphl$BN$Y);
  endspecify
endmodule // NAND2XBX6MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2XBX4MA10TR (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nand (Y, A, Bx);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$BN$Y = 1.0,
      tphl$BN$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (BN *> Y) = (tplh$BN$Y, tphl$BN$Y);
  endspecify
endmodule // NAND2XBX4MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2XBX3MA10TR (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nand (Y, A, Bx);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$BN$Y = 1.0,
      tphl$BN$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (BN *> Y) = (tplh$BN$Y, tphl$BN$Y);
  endspecify
endmodule // NAND2XBX3MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2XBX2MA10TR (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nand (Y, A, Bx);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$BN$Y = 1.0,
      tphl$BN$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (BN *> Y) = (tplh$BN$Y, tphl$BN$Y);
  endspecify
endmodule // NAND2XBX2MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2XBX1P4MA10TR (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nand (Y, A, Bx);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$BN$Y = 1.0,
      tphl$BN$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (BN *> Y) = (tplh$BN$Y, tphl$BN$Y);
  endspecify
endmodule // NAND2XBX1P4MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2XBX1MA10TR (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nand (Y, A, Bx);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$BN$Y = 1.0,
      tphl$BN$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (BN *> Y) = (tplh$BN$Y, tphl$BN$Y);
  endspecify
endmodule // NAND2XBX1MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2XBX0P7MA10TR (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nand (Y, A, Bx);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$BN$Y = 1.0,
      tphl$BN$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (BN *> Y) = (tplh$BN$Y, tphl$BN$Y);
  endspecify
endmodule // NAND2XBX0P7MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2XBX0P5MA10TR (Y, A, BN);
output Y;
input A, BN;

  not (Bx, BN);
  nand (Y, A, Bx);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$BN$Y = 1.0,
      tphl$BN$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (BN *> Y) = (tplh$BN$Y, tphl$BN$Y);
  endspecify
endmodule // NAND2XBX0P5MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2BX8MA10TR (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nand (Y, Ax, B);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2BX8MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2BX6MA10TR (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nand (Y, Ax, B);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2BX6MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2BX4MA10TR (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nand (Y, Ax, B);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2BX4MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2BX3MA10TR (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nand (Y, Ax, B);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2BX3MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2BX2MA10TR (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nand (Y, Ax, B);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2BX2MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2BX1P4MA10TR (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nand (Y, Ax, B);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2BX1P4MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2BX1MA10TR (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nand (Y, Ax, B);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2BX1MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2BX0P7MA10TR (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nand (Y, Ax, B);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2BX0P7MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2BX0P5MA10TR (Y, AN, B);
output Y;
input AN, B;

  not (Ax, AN);
  nand (Y, Ax, B);
  specify
    // delay parameters
    specparam
      tplh$AN$Y = 1.0,
      tphl$AN$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (AN *> Y) = (tplh$AN$Y, tphl$AN$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2BX0P5MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2X8MA10TR (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2X8MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2X8BA10TR (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2X8BA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2X8AA10TR (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2X8AA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2X6MA10TR (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2X6MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2X6BA10TR (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2X6BA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2X6AA10TR (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2X6AA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2X4MA10TR (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2X4MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2X4BA10TR (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2X4BA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2X4AA10TR (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2X4AA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2X3MA10TR (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2X3MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2X3BA10TR (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2X3BA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2X3AA10TR (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2X3AA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2X2MA10TR (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2X2MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2X2BA10TR (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2X2BA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2X2AA10TR (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2X2AA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2X1P4MA10TR (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2X1P4MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2X1P4BA10TR (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2X1P4BA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2X1P4AA10TR (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2X1P4AA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2X1MA10TR (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2X1MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2X1BA10TR (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2X1BA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2X1AA10TR (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2X1AA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2X0P7MA10TR (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2X0P7MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2X0P7BA10TR (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2X0P7BA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2X0P7AA10TR (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2X0P7AA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2X0P5MA10TR (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2X0P5MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2X0P5BA10TR (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2X0P5BA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module NAND2X0P5AA10TR (Y, A, B);
output Y;
input A, B;

  nand (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // NAND2X0P5AA10TR
`endcelldefine
//$Id: mux.genpp,v 1.10 2006/06/19 10:38:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MXT4X3MA10TR (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(Y, A, B, C, D, S0, S1);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0,
      tplh$S1$Y = 1.0,
      tphl$S1$Y = 1.0;
    // path delays
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b0 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b1 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b1 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b0 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b0 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b0 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b1 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b1 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y);
  endspecify

endmodule // MXT4X3MA10TR
`endcelldefine
//$Id: mux.genpp,v 1.10 2006/06/19 10:38:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MXT4X2MA10TR (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(Y, A, B, C, D, S0, S1);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0,
      tplh$S1$Y = 1.0,
      tphl$S1$Y = 1.0;
    // path delays
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b0 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b1 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b1 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b0 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b0 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b0 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b1 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b1 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y);
  endspecify

endmodule // MXT4X2MA10TR
`endcelldefine
//$Id: mux.genpp,v 1.10 2006/06/19 10:38:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MXT4X1P4MA10TR (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(Y, A, B, C, D, S0, S1);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0,
      tplh$S1$Y = 1.0,
      tphl$S1$Y = 1.0;
    // path delays
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b0 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b1 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b1 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b0 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b0 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b0 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b1 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b1 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y);
  endspecify

endmodule // MXT4X1P4MA10TR
`endcelldefine
//$Id: mux.genpp,v 1.10 2006/06/19 10:38:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MXT4X1MA10TR (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(Y, A, B, C, D, S0, S1);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0,
      tplh$S1$Y = 1.0,
      tphl$S1$Y = 1.0;
    // path delays
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b0 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b1 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b1 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b0 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b0 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b0 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b1 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b1 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y);
  endspecify

endmodule // MXT4X1MA10TR
`endcelldefine
//$Id: mux.genpp,v 1.10 2006/06/19 10:38:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MXT4X0P7MA10TR (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(Y, A, B, C, D, S0, S1);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0,
      tplh$S1$Y = 1.0,
      tphl$S1$Y = 1.0;
    // path delays
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b0 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b1 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b1 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b0 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b0 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b0 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b1 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b1 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y);
  endspecify

endmodule // MXT4X0P7MA10TR
`endcelldefine
//$Id: mux.genpp,v 1.10 2006/06/19 10:38:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MXT4X0P5MA10TR (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(Y, A, B, C, D, S0, S1);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0,
      tplh$S1$Y = 1.0,
      tphl$S1$Y = 1.0;
    // path delays
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b0 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b1 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b1 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b0 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b0 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b0 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b1 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b1 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y);
  endspecify

endmodule // MXT4X0P5MA10TR
`endcelldefine
//$Id: mux.genpp,v 1.10 2006/06/19 10:38:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MXT2X6MA10TR (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MXT2X6MA10TR
`endcelldefine
//$Id: mux.genpp,v 1.10 2006/06/19 10:38:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MXT2X4MA10TR (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MXT2X4MA10TR
`endcelldefine
//$Id: mux.genpp,v 1.10 2006/06/19 10:38:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MXT2X3MA10TR (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MXT2X3MA10TR
`endcelldefine
//$Id: mux.genpp,v 1.10 2006/06/19 10:38:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MXT2X2MA10TR (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MXT2X2MA10TR
`endcelldefine
//$Id: mux.genpp,v 1.10 2006/06/19 10:38:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MXT2X1P4MA10TR (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MXT2X1P4MA10TR
`endcelldefine
//$Id: mux.genpp,v 1.10 2006/06/19 10:38:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MXT2X1MA10TR (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MXT2X1MA10TR
`endcelldefine
//$Id: mux.genpp,v 1.10 2006/06/19 10:38:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MXT2X0P7MA10TR (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MXT2X0P7MA10TR
`endcelldefine
//$Id: mux.genpp,v 1.10 2006/06/19 10:38:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MXT2X0P5MA10TR (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MXT2X0P5MA10TR
`endcelldefine
//$Id: mux.genpp,v 1.10 2006/06/19 10:38:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MXIT4X3MA10TR (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      u1(Y, YN);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0,
      tplh$S1$Y = 1.0,
      tphl$S1$Y = 1.0;
    // path delays
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b0 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b1 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b1 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b0 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b0 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b0 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b1 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b1 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y);
  endspecify

endmodule // MXIT4X3MA10TR
`endcelldefine
//$Id: mux.genpp,v 1.10 2006/06/19 10:38:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MXIT4X2MA10TR (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      u1(Y, YN);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0,
      tplh$S1$Y = 1.0,
      tphl$S1$Y = 1.0;
    // path delays
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b0 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b1 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b1 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b0 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b0 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b0 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b1 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b1 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y);
  endspecify

endmodule // MXIT4X2MA10TR
`endcelldefine
//$Id: mux.genpp,v 1.10 2006/06/19 10:38:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MXIT4X1P4MA10TR (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      u1(Y, YN);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0,
      tplh$S1$Y = 1.0,
      tphl$S1$Y = 1.0;
    // path delays
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b0 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b1 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b1 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b0 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b0 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b0 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b1 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b1 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y);
  endspecify

endmodule // MXIT4X1P4MA10TR
`endcelldefine
//$Id: mux.genpp,v 1.10 2006/06/19 10:38:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MXIT4X1MA10TR (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      u1(Y, YN);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0,
      tplh$S1$Y = 1.0,
      tphl$S1$Y = 1.0;
    // path delays
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b0 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b1 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b1 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b0 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b0 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b0 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b1 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b1 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y);
  endspecify

endmodule // MXIT4X1MA10TR
`endcelldefine
//$Id: mux.genpp,v 1.10 2006/06/19 10:38:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MXIT4X0P7MA10TR (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      u1(Y, YN);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0,
      tplh$S1$Y = 1.0,
      tphl$S1$Y = 1.0;
    // path delays
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b0 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b1 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b1 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b0 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b0 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b0 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b1 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b1 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y);
  endspecify

endmodule // MXIT4X0P7MA10TR
`endcelldefine
//$Id: mux.genpp,v 1.10 2006/06/19 10:38:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MXIT4X0P5MA10TR (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;

  udp_mux4 u0(YN, A, B, C, D, S0, S1);
  not      u1(Y, YN);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0,
      tplh$S1$Y = 1.0,
      tphl$S1$Y = 1.0;
    // path delays
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b0 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b0 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b0 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && A == 1'b0 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b1 && S1 == 1'b0 && D == 1'b1 && C == 1'b1 && A == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b0 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b1 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b0 && A == 1'b0 && B == 1'b1 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b0 && S1 == 1'b1 && D == 1'b1 && A == 1'b1 && B == 1'b0 )
       (C *> Y) = (tplh$C$Y, tphl$C$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b0 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b1 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b1 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b0 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b0 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b0 && C == 1'b0 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b1 && B == 1'b0 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S0 == 1'b1 && S1 == 1'b1 && A == 1'b1 && C == 1'b1 && B == 1'b1 )
       (D *> Y) = (tplh$D$Y, tphl$D$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S1 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S0 *> Y) = (tplh$S0$Y, tphl$S0$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b1 && C == 1'b0 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b1 && C == 1'b1 && B == 1'b0 && A == 1'b0 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b0 && D == 1'b0 && C == 1'b0 && B == 1'b0 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y); 
    if (S0 == 1'b1 && D == 1'b0 && C == 1'b1 && B == 1'b1 && A == 1'b1 )
       (S1 *> Y) = (tplh$S1$Y, tphl$S1$Y);
  endspecify

endmodule // MXIT4X0P5MA10TR
`endcelldefine
//$Id: mux.genpp,v 1.10 2006/06/19 10:38:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MXIT2X4MA10TR (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(Y, YN);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MXIT2X4MA10TR
`endcelldefine
//$Id: mux.genpp,v 1.10 2006/06/19 10:38:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MXIT2X3MA10TR (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(Y, YN);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MXIT2X3MA10TR
`endcelldefine
//$Id: mux.genpp,v 1.10 2006/06/19 10:38:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MXIT2X2MA10TR (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(Y, YN);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MXIT2X2MA10TR
`endcelldefine
//$Id: mux.genpp,v 1.10 2006/06/19 10:38:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MXIT2X1P4MA10TR (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(Y, YN);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MXIT2X1P4MA10TR
`endcelldefine
//$Id: mux.genpp,v 1.10 2006/06/19 10:38:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MXIT2X1MA10TR (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(Y, YN);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MXIT2X1MA10TR
`endcelldefine
//$Id: mux.genpp,v 1.10 2006/06/19 10:38:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MXIT2X0P7MA10TR (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(Y, YN);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MXIT2X0P7MA10TR
`endcelldefine
//$Id: mux.genpp,v 1.10 2006/06/19 10:38:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MXIT2X0P5MA10TR (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(YN, A, B, S0);
  not      u1(Y, YN);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MXIT2X0P5MA10TR
`endcelldefine
//$Id: mux.genpp,v 1.10 2006/06/19 10:38:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MX2X8BA10TR (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MX2X8BA10TR
`endcelldefine
//$Id: mux.genpp,v 1.10 2006/06/19 10:38:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MX2X6MA10TR (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MX2X6MA10TR
`endcelldefine
//$Id: mux.genpp,v 1.10 2006/06/19 10:38:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MX2X6BA10TR (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MX2X6BA10TR
`endcelldefine
//$Id: mux.genpp,v 1.10 2006/06/19 10:38:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MX2X4MA10TR (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MX2X4MA10TR
`endcelldefine
//$Id: mux.genpp,v 1.10 2006/06/19 10:38:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MX2X4BA10TR (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MX2X4BA10TR
`endcelldefine
//$Id: mux.genpp,v 1.10 2006/06/19 10:38:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MX2X3MA10TR (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MX2X3MA10TR
`endcelldefine
//$Id: mux.genpp,v 1.10 2006/06/19 10:38:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MX2X3BA10TR (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MX2X3BA10TR
`endcelldefine
//$Id: mux.genpp,v 1.10 2006/06/19 10:38:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MX2X2MA10TR (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MX2X2MA10TR
`endcelldefine
//$Id: mux.genpp,v 1.10 2006/06/19 10:38:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MX2X2BA10TR (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MX2X2BA10TR
`endcelldefine
//$Id: mux.genpp,v 1.10 2006/06/19 10:38:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MX2X1P4MA10TR (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MX2X1P4MA10TR
`endcelldefine
//$Id: mux.genpp,v 1.10 2006/06/19 10:38:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MX2X1P4BA10TR (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MX2X1P4BA10TR
`endcelldefine
//$Id: mux.genpp,v 1.10 2006/06/19 10:38:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MX2X1MA10TR (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MX2X1MA10TR
`endcelldefine
//$Id: mux.genpp,v 1.10 2006/06/19 10:38:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MX2X1BA10TR (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MX2X1BA10TR
`endcelldefine
//$Id: mux.genpp,v 1.10 2006/06/19 10:38:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MX2X0P7MA10TR (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MX2X0P7MA10TR
`endcelldefine
//$Id: mux.genpp,v 1.10 2006/06/19 10:38:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MX2X0P7BA10TR (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MX2X0P7BA10TR
`endcelldefine
//$Id: mux.genpp,v 1.10 2006/06/19 10:38:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MX2X0P5MA10TR (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MX2X0P5MA10TR
`endcelldefine
//$Id: mux.genpp,v 1.10 2006/06/19 10:38:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module MX2X0P5BA10TR (Y, A, B, S0);
output Y;
input A, B, S0;

  udp_mux2 u0(Y, A, B, S0);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$S0$Y = 1.0,
      tphl$S0$Y = 1.0;
    // path delays
     if ((A == 1'b1) && (B == 1'b0))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
     if ((A == 1'b0) && (B == 1'b1))
	(S0 *> Y) = (tplh$S0$Y, tphl$S0$Y);
    if (B == 1'b0 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (B == 1'b1 && S0 == 1'b0 )
       (A *> Y) = (tplh$A$Y, tphl$A$Y); 
    if (A == 1'b0 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y); 
    if (A == 1'b1 && S0 == 1'b1 )
       (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify

endmodule // MX2X0P5BA10TR
`endcelldefine
//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module M2SDFFQNX3MA10TR (QN, D0, D1, S0, SI, SE, CK);
output QN;
input D0, D1, S0, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_mux I0 (nm, D0, D1, S0);
  udp_dff I1 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I2 (n1, nm, SI, SE);
  not     I3 (QN, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  not     I7 (nsel, S0);
  and     I8 (SandRandSEb0, SandR, SEb, nsel);
  and     I9 (SandRandSEb1, SandR, SEb, S0);
  xor     I10 (flag0, nm, SI);
  xor     I12 (D0xorD1, D0, D1);
  and     I13 (flag1, D0xorD1, SandR,SEb);
  specify
    specparam 
      tplh$CK$QN = 1.0,
      tphl$CK$QN = 1.0,
      tsetup$D0$CK = 1.0,
      thold$D0$CK = 0.5,
      tsetup$D1$CK = 1.0,
      thold$D1$CK = 0.5,
      tsetup$S0$CK = 1.0,
      thold$S0$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb0 )
      (posedge CK *> (QN    -: D0)) = (tplh$CK$QN,    tphl$CK$QN);
    if ( SandRandSEb1 )
      (posedge CK *> (QN    -: D1)) = (tplh$CK$QN,    tphl$CK$QN);
    if ( SandRandSE )
      (posedge CK *> (QN    -: SI)) = (tplh$CK$QN,    tphl$CK$QN);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb0 == 1), posedge D0, tsetup$D0$CK  ,thold$D0$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb0 == 1), negedge D0, tsetup$D0$CK  ,thold$D0$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb1 == 1), posedge D1, tsetup$D1$CK  ,thold$D1$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb1 == 1), negedge D1, tsetup$D1$CK  ,thold$D1$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (flag0 == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (flag0 == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (flag1 == 1), posedge S0, tsetup$S0$CK, thold$S0$CK , NOTIFIER);
    $setuphold(posedge CK &&& (flag1 == 1), negedge S0, tsetup$S0$CK, thold$S0$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // M2SDFFQNX3MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module M2SDFFQNX2MA10TR (QN, D0, D1, S0, SI, SE, CK);
output QN;
input D0, D1, S0, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_mux I0 (nm, D0, D1, S0);
  udp_dff I1 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I2 (n1, nm, SI, SE);
  not     I3 (QN, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  not     I7 (nsel, S0);
  and     I8 (SandRandSEb0, SandR, SEb, nsel);
  and     I9 (SandRandSEb1, SandR, SEb, S0);
  xor     I10 (flag0, nm, SI);
  xor     I12 (D0xorD1, D0, D1);
  and     I13 (flag1, D0xorD1, SandR,SEb);
  specify
    specparam 
      tplh$CK$QN = 1.0,
      tphl$CK$QN = 1.0,
      tsetup$D0$CK = 1.0,
      thold$D0$CK = 0.5,
      tsetup$D1$CK = 1.0,
      thold$D1$CK = 0.5,
      tsetup$S0$CK = 1.0,
      thold$S0$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb0 )
      (posedge CK *> (QN    -: D0)) = (tplh$CK$QN,    tphl$CK$QN);
    if ( SandRandSEb1 )
      (posedge CK *> (QN    -: D1)) = (tplh$CK$QN,    tphl$CK$QN);
    if ( SandRandSE )
      (posedge CK *> (QN    -: SI)) = (tplh$CK$QN,    tphl$CK$QN);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb0 == 1), posedge D0, tsetup$D0$CK  ,thold$D0$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb0 == 1), negedge D0, tsetup$D0$CK  ,thold$D0$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb1 == 1), posedge D1, tsetup$D1$CK  ,thold$D1$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb1 == 1), negedge D1, tsetup$D1$CK  ,thold$D1$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (flag0 == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (flag0 == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (flag1 == 1), posedge S0, tsetup$S0$CK, thold$S0$CK , NOTIFIER);
    $setuphold(posedge CK &&& (flag1 == 1), negedge S0, tsetup$S0$CK, thold$S0$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // M2SDFFQNX2MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module M2SDFFQNX1MA10TR (QN, D0, D1, S0, SI, SE, CK);
output QN;
input D0, D1, S0, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_mux I0 (nm, D0, D1, S0);
  udp_dff I1 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I2 (n1, nm, SI, SE);
  not     I3 (QN, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  not     I7 (nsel, S0);
  and     I8 (SandRandSEb0, SandR, SEb, nsel);
  and     I9 (SandRandSEb1, SandR, SEb, S0);
  xor     I10 (flag0, nm, SI);
  xor     I12 (D0xorD1, D0, D1);
  and     I13 (flag1, D0xorD1, SandR,SEb);
  specify
    specparam 
      tplh$CK$QN = 1.0,
      tphl$CK$QN = 1.0,
      tsetup$D0$CK = 1.0,
      thold$D0$CK = 0.5,
      tsetup$D1$CK = 1.0,
      thold$D1$CK = 0.5,
      tsetup$S0$CK = 1.0,
      thold$S0$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb0 )
      (posedge CK *> (QN    -: D0)) = (tplh$CK$QN,    tphl$CK$QN);
    if ( SandRandSEb1 )
      (posedge CK *> (QN    -: D1)) = (tplh$CK$QN,    tphl$CK$QN);
    if ( SandRandSE )
      (posedge CK *> (QN    -: SI)) = (tplh$CK$QN,    tphl$CK$QN);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb0 == 1), posedge D0, tsetup$D0$CK  ,thold$D0$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb0 == 1), negedge D0, tsetup$D0$CK  ,thold$D0$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb1 == 1), posedge D1, tsetup$D1$CK  ,thold$D1$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb1 == 1), negedge D1, tsetup$D1$CK  ,thold$D1$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (flag0 == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (flag0 == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (flag1 == 1), posedge S0, tsetup$S0$CK, thold$S0$CK , NOTIFIER);
    $setuphold(posedge CK &&& (flag1 == 1), negedge S0, tsetup$S0$CK, thold$S0$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // M2SDFFQNX1MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module M2SDFFQNX0P5MA10TR (QN, D0, D1, S0, SI, SE, CK);
output QN;
input D0, D1, S0, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_mux I0 (nm, D0, D1, S0);
  udp_dff I1 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I2 (n1, nm, SI, SE);
  not     I3 (QN, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  not     I7 (nsel, S0);
  and     I8 (SandRandSEb0, SandR, SEb, nsel);
  and     I9 (SandRandSEb1, SandR, SEb, S0);
  xor     I10 (flag0, nm, SI);
  xor     I12 (D0xorD1, D0, D1);
  and     I13 (flag1, D0xorD1, SandR,SEb);
  specify
    specparam 
      tplh$CK$QN = 1.0,
      tphl$CK$QN = 1.0,
      tsetup$D0$CK = 1.0,
      thold$D0$CK = 0.5,
      tsetup$D1$CK = 1.0,
      thold$D1$CK = 0.5,
      tsetup$S0$CK = 1.0,
      thold$S0$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb0 )
      (posedge CK *> (QN    -: D0)) = (tplh$CK$QN,    tphl$CK$QN);
    if ( SandRandSEb1 )
      (posedge CK *> (QN    -: D1)) = (tplh$CK$QN,    tphl$CK$QN);
    if ( SandRandSE )
      (posedge CK *> (QN    -: SI)) = (tplh$CK$QN,    tphl$CK$QN);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb0 == 1), posedge D0, tsetup$D0$CK  ,thold$D0$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb0 == 1), negedge D0, tsetup$D0$CK  ,thold$D0$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb1 == 1), posedge D1, tsetup$D1$CK  ,thold$D1$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb1 == 1), negedge D1, tsetup$D1$CK  ,thold$D1$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (flag0 == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (flag0 == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (flag1 == 1), posedge S0, tsetup$S0$CK, thold$S0$CK , NOTIFIER);
    $setuphold(posedge CK &&& (flag1 == 1), negedge S0, tsetup$S0$CK, thold$S0$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // M2SDFFQNX0P5MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module M2SDFFQX4MA10TR (Q, D0, D1, S0, SI, SE, CK);
output Q;
input D0, D1, S0, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_mux I0 (nm, D0, D1, S0);
  udp_dff I1 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I2 (n1, nm, SI, SE);
  buf     I3 (Q, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  not     I7 (nsel, S0);
  and     I8 (SandRandSEb0, SandR, SEb, nsel);
  and     I9 (SandRandSEb1, SandR, SEb, S0);
  xor     I10 (flag0, nm, SI);
  xor     I12 (D0xorD1, D0, D1);
  and     I13 (flag1, D0xorD1, SandR,SEb);
  specify
    specparam 
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D0$CK = 1.0,
      thold$D0$CK = 0.5,
      tsetup$D1$CK = 1.0,
      thold$D1$CK = 0.5,
      tsetup$S0$CK = 1.0,
      thold$S0$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb0 )
      (posedge CK *> (Q    +: D0)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSEb1 )
      (posedge CK *> (Q    +: D1)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb0 == 1), posedge D0, tsetup$D0$CK  ,thold$D0$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb0 == 1), negedge D0, tsetup$D0$CK  ,thold$D0$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb1 == 1), posedge D1, tsetup$D1$CK  ,thold$D1$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb1 == 1), negedge D1, tsetup$D1$CK  ,thold$D1$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (flag0 == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (flag0 == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (flag1 == 1), posedge S0, tsetup$S0$CK, thold$S0$CK , NOTIFIER);
    $setuphold(posedge CK &&& (flag1 == 1), negedge S0, tsetup$S0$CK, thold$S0$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // M2SDFFQX4MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module M2SDFFQX3MA10TR (Q, D0, D1, S0, SI, SE, CK);
output Q;
input D0, D1, S0, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_mux I0 (nm, D0, D1, S0);
  udp_dff I1 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I2 (n1, nm, SI, SE);
  buf     I3 (Q, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  not     I7 (nsel, S0);
  and     I8 (SandRandSEb0, SandR, SEb, nsel);
  and     I9 (SandRandSEb1, SandR, SEb, S0);
  xor     I10 (flag0, nm, SI);
  xor     I12 (D0xorD1, D0, D1);
  and     I13 (flag1, D0xorD1, SandR,SEb);
  specify
    specparam 
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D0$CK = 1.0,
      thold$D0$CK = 0.5,
      tsetup$D1$CK = 1.0,
      thold$D1$CK = 0.5,
      tsetup$S0$CK = 1.0,
      thold$S0$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb0 )
      (posedge CK *> (Q    +: D0)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSEb1 )
      (posedge CK *> (Q    +: D1)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb0 == 1), posedge D0, tsetup$D0$CK  ,thold$D0$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb0 == 1), negedge D0, tsetup$D0$CK  ,thold$D0$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb1 == 1), posedge D1, tsetup$D1$CK  ,thold$D1$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb1 == 1), negedge D1, tsetup$D1$CK  ,thold$D1$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (flag0 == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (flag0 == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (flag1 == 1), posedge S0, tsetup$S0$CK, thold$S0$CK , NOTIFIER);
    $setuphold(posedge CK &&& (flag1 == 1), negedge S0, tsetup$S0$CK, thold$S0$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // M2SDFFQX3MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module M2SDFFQX2MA10TR (Q, D0, D1, S0, SI, SE, CK);
output Q;
input D0, D1, S0, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_mux I0 (nm, D0, D1, S0);
  udp_dff I1 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I2 (n1, nm, SI, SE);
  buf     I3 (Q, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  not     I7 (nsel, S0);
  and     I8 (SandRandSEb0, SandR, SEb, nsel);
  and     I9 (SandRandSEb1, SandR, SEb, S0);
  xor     I10 (flag0, nm, SI);
  xor     I12 (D0xorD1, D0, D1);
  and     I13 (flag1, D0xorD1, SandR,SEb);
  specify
    specparam 
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D0$CK = 1.0,
      thold$D0$CK = 0.5,
      tsetup$D1$CK = 1.0,
      thold$D1$CK = 0.5,
      tsetup$S0$CK = 1.0,
      thold$S0$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb0 )
      (posedge CK *> (Q    +: D0)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSEb1 )
      (posedge CK *> (Q    +: D1)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb0 == 1), posedge D0, tsetup$D0$CK  ,thold$D0$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb0 == 1), negedge D0, tsetup$D0$CK  ,thold$D0$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb1 == 1), posedge D1, tsetup$D1$CK  ,thold$D1$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb1 == 1), negedge D1, tsetup$D1$CK  ,thold$D1$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (flag0 == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (flag0 == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (flag1 == 1), posedge S0, tsetup$S0$CK, thold$S0$CK , NOTIFIER);
    $setuphold(posedge CK &&& (flag1 == 1), negedge S0, tsetup$S0$CK, thold$S0$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // M2SDFFQX2MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module M2SDFFQX1MA10TR (Q, D0, D1, S0, SI, SE, CK);
output Q;
input D0, D1, S0, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_mux I0 (nm, D0, D1, S0);
  udp_dff I1 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I2 (n1, nm, SI, SE);
  buf     I3 (Q, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  not     I7 (nsel, S0);
  and     I8 (SandRandSEb0, SandR, SEb, nsel);
  and     I9 (SandRandSEb1, SandR, SEb, S0);
  xor     I10 (flag0, nm, SI);
  xor     I12 (D0xorD1, D0, D1);
  and     I13 (flag1, D0xorD1, SandR,SEb);
  specify
    specparam 
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D0$CK = 1.0,
      thold$D0$CK = 0.5,
      tsetup$D1$CK = 1.0,
      thold$D1$CK = 0.5,
      tsetup$S0$CK = 1.0,
      thold$S0$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb0 )
      (posedge CK *> (Q    +: D0)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSEb1 )
      (posedge CK *> (Q    +: D1)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb0 == 1), posedge D0, tsetup$D0$CK  ,thold$D0$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb0 == 1), negedge D0, tsetup$D0$CK  ,thold$D0$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb1 == 1), posedge D1, tsetup$D1$CK  ,thold$D1$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb1 == 1), negedge D1, tsetup$D1$CK  ,thold$D1$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (flag0 == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (flag0 == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (flag1 == 1), posedge S0, tsetup$S0$CK, thold$S0$CK , NOTIFIER);
    $setuphold(posedge CK &&& (flag1 == 1), negedge S0, tsetup$S0$CK, thold$S0$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // M2SDFFQX1MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module M2SDFFQX0P5MA10TR (Q, D0, D1, S0, SI, SE, CK);
output Q;
input D0, D1, S0, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  udp_mux I0 (nm, D0, D1, S0);
  udp_dff I1 (n0, n1, clk, xRN, xSN, NOTIFIER);
  udp_mux I2 (n1, nm, SI, SE);
  buf     I3 (Q, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  not     I7 (nsel, S0);
  and     I8 (SandRandSEb0, SandR, SEb, nsel);
  and     I9 (SandRandSEb1, SandR, SEb, S0);
  xor     I10 (flag0, nm, SI);
  xor     I12 (D0xorD1, D0, D1);
  and     I13 (flag1, D0xorD1, SandR,SEb);
  specify
    specparam 
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$D0$CK = 1.0,
      thold$D0$CK = 0.5,
      tsetup$D1$CK = 1.0,
      thold$D1$CK = 0.5,
      tsetup$S0$CK = 1.0,
      thold$S0$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEb0 )
      (posedge CK *> (Q    +: D0)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSEb1 )
      (posedge CK *> (Q    +: D1)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb0 == 1), posedge D0, tsetup$D0$CK  ,thold$D0$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb0 == 1), negedge D0, tsetup$D0$CK  ,thold$D0$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb1 == 1), posedge D1, tsetup$D1$CK  ,thold$D1$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb1 == 1), negedge D1, tsetup$D1$CK  ,thold$D1$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (flag0 == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (flag0 == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (flag1 == 1), posedge S0, tsetup$S0$CK, thold$S0$CK , NOTIFIER);
    $setuphold(posedge CK &&& (flag1 == 1), negedge S0, tsetup$S0$CK, thold$S0$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // M2SDFFQX0P5MA10TR
`endcelldefine
	

//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module M2DFFQNX3MA10TR (QN, D0, D1, S0, CK);
output QN;
input  D0, D1, S0, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_mux2 I0 (nm, D0, D1, S0);
  udp_dff  I1 (n0, nm, clk, xRN, xSN, NOTIFIER);
  not      I5 (QN, n0);
  not      I2 (nsel,S0);
  and      I3 (flag0, xRN, xSN, nsel);
  and      I4 (flag1, xRN, xSN, S0);
  xor      I6 (D0xorD1, D0, D1);
  and      I7 (flag, D0xorD1, xRN, xSN);
  and      I8 (SandR,xRN, xSN);
  specify
    specparam
    tplh$CK$QN	= 1.0,
    tphl$CK$QN	= 1.0,
    tsetup$D0$CK	= 1.0,
    thold$D0$CK	= 0.5,
    tsetup$D1$CK	= 1.0,
    thold$D1$CK	= 0.5,
    tsetup$S0$CK	= 1.0,
    thold$S0$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;

    if (flag0)
      (posedge CK *> (QN -: D0)) = (tplh$CK$QN,    tphl$CK$QN);
    if (flag1)
      (posedge CK *> (QN -: D1)) = (tplh$CK$QN,    tphl$CK$QN);

    $setuphold(posedge CK &&& (flag0 == 1), posedge D0, tsetup$D0$CK, thold$D0$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag0 == 1), negedge D0, tsetup$D0$CK, thold$D0$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag1 == 1), posedge D1, tsetup$D1$CK, thold$D1$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag1 == 1), negedge D1, tsetup$D1$CK, thold$D1$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), posedge S0, tsetup$S0$CK, thold$S0$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge S0, tsetup$S0$CK, thold$S0$CK, NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // M2DFFQNX3MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module M2DFFQNX2MA10TR (QN, D0, D1, S0, CK);
output QN;
input  D0, D1, S0, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_mux2 I0 (nm, D0, D1, S0);
  udp_dff  I1 (n0, nm, clk, xRN, xSN, NOTIFIER);
  not      I5 (QN, n0);
  not      I2 (nsel,S0);
  and      I3 (flag0, xRN, xSN, nsel);
  and      I4 (flag1, xRN, xSN, S0);
  xor      I6 (D0xorD1, D0, D1);
  and      I7 (flag, D0xorD1, xRN, xSN);
  and      I8 (SandR,xRN, xSN);
  specify
    specparam
    tplh$CK$QN	= 1.0,
    tphl$CK$QN	= 1.0,
    tsetup$D0$CK	= 1.0,
    thold$D0$CK	= 0.5,
    tsetup$D1$CK	= 1.0,
    thold$D1$CK	= 0.5,
    tsetup$S0$CK	= 1.0,
    thold$S0$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;

    if (flag0)
      (posedge CK *> (QN -: D0)) = (tplh$CK$QN,    tphl$CK$QN);
    if (flag1)
      (posedge CK *> (QN -: D1)) = (tplh$CK$QN,    tphl$CK$QN);

    $setuphold(posedge CK &&& (flag0 == 1), posedge D0, tsetup$D0$CK, thold$D0$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag0 == 1), negedge D0, tsetup$D0$CK, thold$D0$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag1 == 1), posedge D1, tsetup$D1$CK, thold$D1$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag1 == 1), negedge D1, tsetup$D1$CK, thold$D1$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), posedge S0, tsetup$S0$CK, thold$S0$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge S0, tsetup$S0$CK, thold$S0$CK, NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // M2DFFQNX2MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module M2DFFQNX1MA10TR (QN, D0, D1, S0, CK);
output QN;
input  D0, D1, S0, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_mux2 I0 (nm, D0, D1, S0);
  udp_dff  I1 (n0, nm, clk, xRN, xSN, NOTIFIER);
  not      I5 (QN, n0);
  not      I2 (nsel,S0);
  and      I3 (flag0, xRN, xSN, nsel);
  and      I4 (flag1, xRN, xSN, S0);
  xor      I6 (D0xorD1, D0, D1);
  and      I7 (flag, D0xorD1, xRN, xSN);
  and      I8 (SandR,xRN, xSN);
  specify
    specparam
    tplh$CK$QN	= 1.0,
    tphl$CK$QN	= 1.0,
    tsetup$D0$CK	= 1.0,
    thold$D0$CK	= 0.5,
    tsetup$D1$CK	= 1.0,
    thold$D1$CK	= 0.5,
    tsetup$S0$CK	= 1.0,
    thold$S0$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;

    if (flag0)
      (posedge CK *> (QN -: D0)) = (tplh$CK$QN,    tphl$CK$QN);
    if (flag1)
      (posedge CK *> (QN -: D1)) = (tplh$CK$QN,    tphl$CK$QN);

    $setuphold(posedge CK &&& (flag0 == 1), posedge D0, tsetup$D0$CK, thold$D0$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag0 == 1), negedge D0, tsetup$D0$CK, thold$D0$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag1 == 1), posedge D1, tsetup$D1$CK, thold$D1$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag1 == 1), negedge D1, tsetup$D1$CK, thold$D1$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), posedge S0, tsetup$S0$CK, thold$S0$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge S0, tsetup$S0$CK, thold$S0$CK, NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // M2DFFQNX1MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module M2DFFQNX0P5MA10TR (QN, D0, D1, S0, CK);
output QN;
input  D0, D1, S0, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_mux2 I0 (nm, D0, D1, S0);
  udp_dff  I1 (n0, nm, clk, xRN, xSN, NOTIFIER);
  not      I5 (QN, n0);
  not      I2 (nsel,S0);
  and      I3 (flag0, xRN, xSN, nsel);
  and      I4 (flag1, xRN, xSN, S0);
  xor      I6 (D0xorD1, D0, D1);
  and      I7 (flag, D0xorD1, xRN, xSN);
  and      I8 (SandR,xRN, xSN);
  specify
    specparam
    tplh$CK$QN	= 1.0,
    tphl$CK$QN	= 1.0,
    tsetup$D0$CK	= 1.0,
    thold$D0$CK	= 0.5,
    tsetup$D1$CK	= 1.0,
    thold$D1$CK	= 0.5,
    tsetup$S0$CK	= 1.0,
    thold$S0$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;

    if (flag0)
      (posedge CK *> (QN -: D0)) = (tplh$CK$QN,    tphl$CK$QN);
    if (flag1)
      (posedge CK *> (QN -: D1)) = (tplh$CK$QN,    tphl$CK$QN);

    $setuphold(posedge CK &&& (flag0 == 1), posedge D0, tsetup$D0$CK, thold$D0$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag0 == 1), negedge D0, tsetup$D0$CK, thold$D0$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag1 == 1), posedge D1, tsetup$D1$CK, thold$D1$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag1 == 1), negedge D1, tsetup$D1$CK, thold$D1$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), posedge S0, tsetup$S0$CK, thold$S0$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge S0, tsetup$S0$CK, thold$S0$CK, NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // M2DFFQNX0P5MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module M2DFFQX4MA10TR (Q, D0, D1, S0, CK);
output Q;
input  D0, D1, S0, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_mux2 I0 (nm, D0, D1, S0);
  udp_dff  I1 (n0, nm, clk, xRN, xSN, NOTIFIER);
  buf      I5 (Q, n0);
  not      I2 (nsel,S0);
  and      I3 (flag0, xRN, xSN, nsel);
  and      I4 (flag1, xRN, xSN, S0);
  xor      I6 (D0xorD1, D0, D1);
  and      I7 (flag, D0xorD1, xRN, xSN);
  and      I8 (SandR,xRN, xSN);
  specify
    specparam
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D0$CK	= 1.0,
    thold$D0$CK	= 0.5,
    tsetup$D1$CK	= 1.0,
    thold$D1$CK	= 0.5,
    tsetup$S0$CK	= 1.0,
    thold$S0$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;

    if (flag0)
      (posedge CK *> (Q +: D0)) = (tplh$CK$Q,    tphl$CK$Q);
    if (flag1)
      (posedge CK *> (Q +: D1)) = (tplh$CK$Q,    tphl$CK$Q);

    $setuphold(posedge CK &&& (flag0 == 1), posedge D0, tsetup$D0$CK, thold$D0$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag0 == 1), negedge D0, tsetup$D0$CK, thold$D0$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag1 == 1), posedge D1, tsetup$D1$CK, thold$D1$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag1 == 1), negedge D1, tsetup$D1$CK, thold$D1$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), posedge S0, tsetup$S0$CK, thold$S0$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge S0, tsetup$S0$CK, thold$S0$CK, NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // M2DFFQX4MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module M2DFFQX3MA10TR (Q, D0, D1, S0, CK);
output Q;
input  D0, D1, S0, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_mux2 I0 (nm, D0, D1, S0);
  udp_dff  I1 (n0, nm, clk, xRN, xSN, NOTIFIER);
  buf      I5 (Q, n0);
  not      I2 (nsel,S0);
  and      I3 (flag0, xRN, xSN, nsel);
  and      I4 (flag1, xRN, xSN, S0);
  xor      I6 (D0xorD1, D0, D1);
  and      I7 (flag, D0xorD1, xRN, xSN);
  and      I8 (SandR,xRN, xSN);
  specify
    specparam
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D0$CK	= 1.0,
    thold$D0$CK	= 0.5,
    tsetup$D1$CK	= 1.0,
    thold$D1$CK	= 0.5,
    tsetup$S0$CK	= 1.0,
    thold$S0$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;

    if (flag0)
      (posedge CK *> (Q +: D0)) = (tplh$CK$Q,    tphl$CK$Q);
    if (flag1)
      (posedge CK *> (Q +: D1)) = (tplh$CK$Q,    tphl$CK$Q);

    $setuphold(posedge CK &&& (flag0 == 1), posedge D0, tsetup$D0$CK, thold$D0$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag0 == 1), negedge D0, tsetup$D0$CK, thold$D0$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag1 == 1), posedge D1, tsetup$D1$CK, thold$D1$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag1 == 1), negedge D1, tsetup$D1$CK, thold$D1$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), posedge S0, tsetup$S0$CK, thold$S0$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge S0, tsetup$S0$CK, thold$S0$CK, NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // M2DFFQX3MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module M2DFFQX2MA10TR (Q, D0, D1, S0, CK);
output Q;
input  D0, D1, S0, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_mux2 I0 (nm, D0, D1, S0);
  udp_dff  I1 (n0, nm, clk, xRN, xSN, NOTIFIER);
  buf      I5 (Q, n0);
  not      I2 (nsel,S0);
  and      I3 (flag0, xRN, xSN, nsel);
  and      I4 (flag1, xRN, xSN, S0);
  xor      I6 (D0xorD1, D0, D1);
  and      I7 (flag, D0xorD1, xRN, xSN);
  and      I8 (SandR,xRN, xSN);
  specify
    specparam
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D0$CK	= 1.0,
    thold$D0$CK	= 0.5,
    tsetup$D1$CK	= 1.0,
    thold$D1$CK	= 0.5,
    tsetup$S0$CK	= 1.0,
    thold$S0$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;

    if (flag0)
      (posedge CK *> (Q +: D0)) = (tplh$CK$Q,    tphl$CK$Q);
    if (flag1)
      (posedge CK *> (Q +: D1)) = (tplh$CK$Q,    tphl$CK$Q);

    $setuphold(posedge CK &&& (flag0 == 1), posedge D0, tsetup$D0$CK, thold$D0$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag0 == 1), negedge D0, tsetup$D0$CK, thold$D0$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag1 == 1), posedge D1, tsetup$D1$CK, thold$D1$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag1 == 1), negedge D1, tsetup$D1$CK, thold$D1$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), posedge S0, tsetup$S0$CK, thold$S0$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge S0, tsetup$S0$CK, thold$S0$CK, NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // M2DFFQX2MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module M2DFFQX1MA10TR (Q, D0, D1, S0, CK);
output Q;
input  D0, D1, S0, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_mux2 I0 (nm, D0, D1, S0);
  udp_dff  I1 (n0, nm, clk, xRN, xSN, NOTIFIER);
  buf      I5 (Q, n0);
  not      I2 (nsel,S0);
  and      I3 (flag0, xRN, xSN, nsel);
  and      I4 (flag1, xRN, xSN, S0);
  xor      I6 (D0xorD1, D0, D1);
  and      I7 (flag, D0xorD1, xRN, xSN);
  and      I8 (SandR,xRN, xSN);
  specify
    specparam
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D0$CK	= 1.0,
    thold$D0$CK	= 0.5,
    tsetup$D1$CK	= 1.0,
    thold$D1$CK	= 0.5,
    tsetup$S0$CK	= 1.0,
    thold$S0$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;

    if (flag0)
      (posedge CK *> (Q +: D0)) = (tplh$CK$Q,    tphl$CK$Q);
    if (flag1)
      (posedge CK *> (Q +: D1)) = (tplh$CK$Q,    tphl$CK$Q);

    $setuphold(posedge CK &&& (flag0 == 1), posedge D0, tsetup$D0$CK, thold$D0$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag0 == 1), negedge D0, tsetup$D0$CK, thold$D0$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag1 == 1), posedge D1, tsetup$D1$CK, thold$D1$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag1 == 1), negedge D1, tsetup$D1$CK, thold$D1$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), posedge S0, tsetup$S0$CK, thold$S0$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge S0, tsetup$S0$CK, thold$S0$CK, NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // M2DFFQX1MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module M2DFFQX0P5MA10TR (Q, D0, D1, S0, CK);
output Q;
input  D0, D1, S0, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_mux2 I0 (nm, D0, D1, S0);
  udp_dff  I1 (n0, nm, clk, xRN, xSN, NOTIFIER);
  buf      I5 (Q, n0);
  not      I2 (nsel,S0);
  and      I3 (flag0, xRN, xSN, nsel);
  and      I4 (flag1, xRN, xSN, S0);
  xor      I6 (D0xorD1, D0, D1);
  and      I7 (flag, D0xorD1, xRN, xSN);
  and      I8 (SandR,xRN, xSN);
  specify
    specparam
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D0$CK	= 1.0,
    thold$D0$CK	= 0.5,
    tsetup$D1$CK	= 1.0,
    thold$D1$CK	= 0.5,
    tsetup$S0$CK	= 1.0,
    thold$S0$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;

    if (flag0)
      (posedge CK *> (Q +: D0)) = (tplh$CK$Q,    tphl$CK$Q);
    if (flag1)
      (posedge CK *> (Q +: D1)) = (tplh$CK$Q,    tphl$CK$Q);

    $setuphold(posedge CK &&& (flag0 == 1), posedge D0, tsetup$D0$CK, thold$D0$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag0 == 1), negedge D0, tsetup$D0$CK, thold$D0$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag1 == 1), posedge D1, tsetup$D1$CK, thold$D1$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag1 == 1), negedge D1, tsetup$D1$CK, thold$D1$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), posedge S0, tsetup$S0$CK, thold$S0$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge S0, tsetup$S0$CK, thold$S0$CK, NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // M2DFFQX0P5MA10TR
`endcelldefine


//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATSQNX4MA10TR (QN, D, G, SN);
output  QN;
input  D, G, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

buf       XX0 (xSN, SN);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
not I3(clk,G);
buf I4(flgclk,G);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$QN   = 1.0,
      tphl$D$QN   = 1.0,
      tplh$G$QN   = 1.0,
      tphl$G$QN   = 1.0,
      tplh$SN$QN   = 1.0,
      tphl$SN$QN   = 1.0,
      tsetup$D$G = 1.0,
      thold$D$G  = 0.5,
      tsetup$D$SN = 1.0,
      thold$D$SN  = 0.5,
      tsetup$G$SN = 1.0,
      thold$G$SN  = 0.5,
      tsetup$SN$G = 1.0,
      thold$SN$G  = 0.5,
      tminpwl$SN = 1.0,
      tminpwh$G  = 1.0,
      tperiod$G  = 1.0;
    // path delays
    if (SandR)
      (posedge G *> (QN    -: D)) = (tplh$G$QN,    tphl$G$QN);
    if (SandRandCLK)
      ( D *> QN ) = (tplh$D$QN, tphl$D$QN );
    $setuphold(negedge G, posedge SN, tsetup$SN$G,thold$SN$G, NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    // timing checks 2
    $setuphold(negedge G &&& (SandR == 1), posedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $setuphold(negedge G &&& (SandR == 1), negedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $width(posedge G &&& (SandR == 1), tminpwh$G, 0, NOTIFIER);
    $period(posedge G &&& (SandR == 1), tperiod$G, NOTIFIER);
    if (D == 1'b0 && G == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN);
    if (D == 1'b0 && G == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN);
    if (D == 1'b1 && G == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN);

   endspecify
endmodule //LATSQNX4MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATSQNX3MA10TR (QN, D, G, SN);
output  QN;
input  D, G, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

buf       XX0 (xSN, SN);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
not I3(clk,G);
buf I4(flgclk,G);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$QN   = 1.0,
      tphl$D$QN   = 1.0,
      tplh$G$QN   = 1.0,
      tphl$G$QN   = 1.0,
      tplh$SN$QN   = 1.0,
      tphl$SN$QN   = 1.0,
      tsetup$D$G = 1.0,
      thold$D$G  = 0.5,
      tsetup$D$SN = 1.0,
      thold$D$SN  = 0.5,
      tsetup$G$SN = 1.0,
      thold$G$SN  = 0.5,
      tsetup$SN$G = 1.0,
      thold$SN$G  = 0.5,
      tminpwl$SN = 1.0,
      tminpwh$G  = 1.0,
      tperiod$G  = 1.0;
    // path delays
    if (SandR)
      (posedge G *> (QN    -: D)) = (tplh$G$QN,    tphl$G$QN);
    if (SandRandCLK)
      ( D *> QN ) = (tplh$D$QN, tphl$D$QN );
    $setuphold(negedge G, posedge SN, tsetup$SN$G,thold$SN$G, NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    // timing checks 2
    $setuphold(negedge G &&& (SandR == 1), posedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $setuphold(negedge G &&& (SandR == 1), negedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $width(posedge G &&& (SandR == 1), tminpwh$G, 0, NOTIFIER);
    $period(posedge G &&& (SandR == 1), tperiod$G, NOTIFIER);
    if (D == 1'b0 && G == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN);
    if (D == 1'b0 && G == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN);
    if (D == 1'b1 && G == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN);

   endspecify
endmodule //LATSQNX3MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATSQNX2MA10TR (QN, D, G, SN);
output  QN;
input  D, G, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

buf       XX0 (xSN, SN);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
not I3(clk,G);
buf I4(flgclk,G);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$QN   = 1.0,
      tphl$D$QN   = 1.0,
      tplh$G$QN   = 1.0,
      tphl$G$QN   = 1.0,
      tplh$SN$QN   = 1.0,
      tphl$SN$QN   = 1.0,
      tsetup$D$G = 1.0,
      thold$D$G  = 0.5,
      tsetup$D$SN = 1.0,
      thold$D$SN  = 0.5,
      tsetup$G$SN = 1.0,
      thold$G$SN  = 0.5,
      tsetup$SN$G = 1.0,
      thold$SN$G  = 0.5,
      tminpwl$SN = 1.0,
      tminpwh$G  = 1.0,
      tperiod$G  = 1.0;
    // path delays
    if (SandR)
      (posedge G *> (QN    -: D)) = (tplh$G$QN,    tphl$G$QN);
    if (SandRandCLK)
      ( D *> QN ) = (tplh$D$QN, tphl$D$QN );
    $setuphold(negedge G, posedge SN, tsetup$SN$G,thold$SN$G, NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    // timing checks 2
    $setuphold(negedge G &&& (SandR == 1), posedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $setuphold(negedge G &&& (SandR == 1), negedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $width(posedge G &&& (SandR == 1), tminpwh$G, 0, NOTIFIER);
    $period(posedge G &&& (SandR == 1), tperiod$G, NOTIFIER);
    if (D == 1'b0 && G == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN);
    if (D == 1'b0 && G == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN);
    if (D == 1'b1 && G == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN);

   endspecify
endmodule //LATSQNX2MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATSQNX1MA10TR (QN, D, G, SN);
output  QN;
input  D, G, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

buf       XX0 (xSN, SN);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
not I3(clk,G);
buf I4(flgclk,G);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$QN   = 1.0,
      tphl$D$QN   = 1.0,
      tplh$G$QN   = 1.0,
      tphl$G$QN   = 1.0,
      tplh$SN$QN   = 1.0,
      tphl$SN$QN   = 1.0,
      tsetup$D$G = 1.0,
      thold$D$G  = 0.5,
      tsetup$D$SN = 1.0,
      thold$D$SN  = 0.5,
      tsetup$G$SN = 1.0,
      thold$G$SN  = 0.5,
      tsetup$SN$G = 1.0,
      thold$SN$G  = 0.5,
      tminpwl$SN = 1.0,
      tminpwh$G  = 1.0,
      tperiod$G  = 1.0;
    // path delays
    if (SandR)
      (posedge G *> (QN    -: D)) = (tplh$G$QN,    tphl$G$QN);
    if (SandRandCLK)
      ( D *> QN ) = (tplh$D$QN, tphl$D$QN );
    $setuphold(negedge G, posedge SN, tsetup$SN$G,thold$SN$G, NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    // timing checks 2
    $setuphold(negedge G &&& (SandR == 1), posedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $setuphold(negedge G &&& (SandR == 1), negedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $width(posedge G &&& (SandR == 1), tminpwh$G, 0, NOTIFIER);
    $period(posedge G &&& (SandR == 1), tperiod$G, NOTIFIER);
    if (D == 1'b0 && G == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN);
    if (D == 1'b0 && G == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN);
    if (D == 1'b1 && G == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN);

   endspecify
endmodule //LATSQNX1MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATSQNX0P5MA10TR (QN, D, G, SN);
output  QN;
input  D, G, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

buf       XX0 (xSN, SN);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
not I3(clk,G);
buf I4(flgclk,G);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$QN   = 1.0,
      tphl$D$QN   = 1.0,
      tplh$G$QN   = 1.0,
      tphl$G$QN   = 1.0,
      tplh$SN$QN   = 1.0,
      tphl$SN$QN   = 1.0,
      tsetup$D$G = 1.0,
      thold$D$G  = 0.5,
      tsetup$D$SN = 1.0,
      thold$D$SN  = 0.5,
      tsetup$G$SN = 1.0,
      thold$G$SN  = 0.5,
      tsetup$SN$G = 1.0,
      thold$SN$G  = 0.5,
      tminpwl$SN = 1.0,
      tminpwh$G  = 1.0,
      tperiod$G  = 1.0;
    // path delays
    if (SandR)
      (posedge G *> (QN    -: D)) = (tplh$G$QN,    tphl$G$QN);
    if (SandRandCLK)
      ( D *> QN ) = (tplh$D$QN, tphl$D$QN );
    $setuphold(negedge G, posedge SN, tsetup$SN$G,thold$SN$G, NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    // timing checks 2
    $setuphold(negedge G &&& (SandR == 1), posedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $setuphold(negedge G &&& (SandR == 1), negedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $width(posedge G &&& (SandR == 1), tminpwh$G, 0, NOTIFIER);
    $period(posedge G &&& (SandR == 1), tperiod$G, NOTIFIER);
    if (D == 1'b0 && G == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN);
    if (D == 1'b0 && G == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN);
    if (D == 1'b1 && G == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN);

   endspecify
endmodule //LATSQNX0P5MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATSPQX3MA10TR (Q, D, G, S);
output  Q;
input  D, G, S;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

not       XX0 (xSN, S);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
not I3(clk,G);
buf I4(flgclk,G);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$Q   = 1.0,
      tphl$D$Q   = 1.0,
      tplh$G$Q   = 1.0,
      tphl$G$Q   = 1.0,
      tplh$S$Q   = 1.0,
      tphl$S$Q   = 1.0,
      tsetup$D$G = 1.0,
      thold$D$G  = 0.5,
      tsetup$D$S = 1.0,
      thold$D$S  = 0.5,
      tsetup$G$S = 1.0,
      thold$G$S  = 0.5,
      tsetup$S$G = 1.0,
      thold$S$G  = 0.5,
      tminpwh$S   = 1.0,
      tminpwh$G  = 1.0,
      tperiod$G  = 1.0;
    // path delays
    if (SandR)
      (posedge G *> (Q    +: D)) = (tplh$G$Q,    tphl$G$Q);
    if (SandRandCLK)
      ( D *> Q ) = (tplh$D$Q, tphl$D$Q );
    $setuphold(negedge G, negedge S, tsetup$S$G,thold$S$G, NOTIFIER);
    $width(posedge S, tminpwh$S, 0, NOTIFIER);
    // timing checks 6
    $setuphold(negedge G &&& (SandR == 1), posedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $setuphold(negedge G &&& (SandR == 1), negedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $width(posedge G &&& (SandR == 1), tminpwh$G, 0, NOTIFIER);
    $period(posedge G &&& (SandR == 1), tperiod$G, NOTIFIER);
    if (D == 1'b0 && G == 1'b0 )
       (posedge  S *> (Q +: 1'b1)) = ( tphl$S$Q);
    if (D == 1'b0 && G == 1'b1 )
       (posedge  S *> (Q +: 1'b1)) = (tplh$S$Q, tphl$S$Q);
    if (D == 1'b1 && G == 1'b0 )
       (posedge  S *> (Q +: 1'b1)) = ( tphl$S$Q);

   endspecify
endmodule //LATSPQX3MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATSPQX2MA10TR (Q, D, G, S);
output  Q;
input  D, G, S;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

not       XX0 (xSN, S);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
not I3(clk,G);
buf I4(flgclk,G);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$Q   = 1.0,
      tphl$D$Q   = 1.0,
      tplh$G$Q   = 1.0,
      tphl$G$Q   = 1.0,
      tplh$S$Q   = 1.0,
      tphl$S$Q   = 1.0,
      tsetup$D$G = 1.0,
      thold$D$G  = 0.5,
      tsetup$D$S = 1.0,
      thold$D$S  = 0.5,
      tsetup$G$S = 1.0,
      thold$G$S  = 0.5,
      tsetup$S$G = 1.0,
      thold$S$G  = 0.5,
      tminpwh$S   = 1.0,
      tminpwh$G  = 1.0,
      tperiod$G  = 1.0;
    // path delays
    if (SandR)
      (posedge G *> (Q    +: D)) = (tplh$G$Q,    tphl$G$Q);
    if (SandRandCLK)
      ( D *> Q ) = (tplh$D$Q, tphl$D$Q );
    $setuphold(negedge G, negedge S, tsetup$S$G,thold$S$G, NOTIFIER);
    $width(posedge S, tminpwh$S, 0, NOTIFIER);
    // timing checks 6
    $setuphold(negedge G &&& (SandR == 1), posedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $setuphold(negedge G &&& (SandR == 1), negedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $width(posedge G &&& (SandR == 1), tminpwh$G, 0, NOTIFIER);
    $period(posedge G &&& (SandR == 1), tperiod$G, NOTIFIER);
    if (D == 1'b0 && G == 1'b0 )
       (posedge  S *> (Q +: 1'b1)) = ( tphl$S$Q);
    if (D == 1'b0 && G == 1'b1 )
       (posedge  S *> (Q +: 1'b1)) = (tplh$S$Q, tphl$S$Q);
    if (D == 1'b1 && G == 1'b0 )
       (posedge  S *> (Q +: 1'b1)) = ( tphl$S$Q);

   endspecify
endmodule //LATSPQX2MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATSPQX1MA10TR (Q, D, G, S);
output  Q;
input  D, G, S;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

not       XX0 (xSN, S);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
not I3(clk,G);
buf I4(flgclk,G);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$Q   = 1.0,
      tphl$D$Q   = 1.0,
      tplh$G$Q   = 1.0,
      tphl$G$Q   = 1.0,
      tplh$S$Q   = 1.0,
      tphl$S$Q   = 1.0,
      tsetup$D$G = 1.0,
      thold$D$G  = 0.5,
      tsetup$D$S = 1.0,
      thold$D$S  = 0.5,
      tsetup$G$S = 1.0,
      thold$G$S  = 0.5,
      tsetup$S$G = 1.0,
      thold$S$G  = 0.5,
      tminpwh$S   = 1.0,
      tminpwh$G  = 1.0,
      tperiod$G  = 1.0;
    // path delays
    if (SandR)
      (posedge G *> (Q    +: D)) = (tplh$G$Q,    tphl$G$Q);
    if (SandRandCLK)
      ( D *> Q ) = (tplh$D$Q, tphl$D$Q );
    $setuphold(negedge G, negedge S, tsetup$S$G,thold$S$G, NOTIFIER);
    $width(posedge S, tminpwh$S, 0, NOTIFIER);
    // timing checks 6
    $setuphold(negedge G &&& (SandR == 1), posedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $setuphold(negedge G &&& (SandR == 1), negedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $width(posedge G &&& (SandR == 1), tminpwh$G, 0, NOTIFIER);
    $period(posedge G &&& (SandR == 1), tperiod$G, NOTIFIER);
    if (D == 1'b0 && G == 1'b0 )
       (posedge  S *> (Q +: 1'b1)) = ( tphl$S$Q);
    if (D == 1'b0 && G == 1'b1 )
       (posedge  S *> (Q +: 1'b1)) = (tplh$S$Q, tphl$S$Q);
    if (D == 1'b1 && G == 1'b0 )
       (posedge  S *> (Q +: 1'b1)) = ( tphl$S$Q);

   endspecify
endmodule //LATSPQX1MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATSPQX0P5MA10TR (Q, D, G, S);
output  Q;
input  D, G, S;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

not       XX0 (xSN, S);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
not I3(clk,G);
buf I4(flgclk,G);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$Q   = 1.0,
      tphl$D$Q   = 1.0,
      tplh$G$Q   = 1.0,
      tphl$G$Q   = 1.0,
      tplh$S$Q   = 1.0,
      tphl$S$Q   = 1.0,
      tsetup$D$G = 1.0,
      thold$D$G  = 0.5,
      tsetup$D$S = 1.0,
      thold$D$S  = 0.5,
      tsetup$G$S = 1.0,
      thold$G$S  = 0.5,
      tsetup$S$G = 1.0,
      thold$S$G  = 0.5,
      tminpwh$S   = 1.0,
      tminpwh$G  = 1.0,
      tperiod$G  = 1.0;
    // path delays
    if (SandR)
      (posedge G *> (Q    +: D)) = (tplh$G$Q,    tphl$G$Q);
    if (SandRandCLK)
      ( D *> Q ) = (tplh$D$Q, tphl$D$Q );
    $setuphold(negedge G, negedge S, tsetup$S$G,thold$S$G, NOTIFIER);
    $width(posedge S, tminpwh$S, 0, NOTIFIER);
    // timing checks 6
    $setuphold(negedge G &&& (SandR == 1), posedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $setuphold(negedge G &&& (SandR == 1), negedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $width(posedge G &&& (SandR == 1), tminpwh$G, 0, NOTIFIER);
    $period(posedge G &&& (SandR == 1), tperiod$G, NOTIFIER);
    if (D == 1'b0 && G == 1'b0 )
       (posedge  S *> (Q +: 1'b1)) = ( tphl$S$Q);
    if (D == 1'b0 && G == 1'b1 )
       (posedge  S *> (Q +: 1'b1)) = (tplh$S$Q, tphl$S$Q);
    if (D == 1'b1 && G == 1'b0 )
       (posedge  S *> (Q +: 1'b1)) = ( tphl$S$Q);

   endspecify
endmodule //LATSPQX0P5MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATRQX3MA10TR (Q, D, G, RN);
output  Q;
input  D, G, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

buf       XX0 (xRN, RN);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
not I3(clk,G);
buf I4(flgclk,G);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$Q   = 1.0,
      tphl$D$Q   = 1.0,
      tplh$G$Q   = 1.0,
      tphl$G$Q   = 1.0,
      tplh$RN$Q   = 1.0,
      tphl$RN$Q   = 1.0,
      tsetup$D$G = 1.0,
      thold$D$G  = 0.5,
      tsetup$D$RN = 1.0,
      thold$D$RN  = 0.5,
      tsetup$G$RN = 1.0,
      thold$G$RN  = 0.5,
      tsetup$RN$G = 1.0,
      thold$RN$G  = 0.5,
      tminpwl$RN    = 1.0,
      tminpwh$G  = 1.0,
      tperiod$G  = 1.0;
    // path delays
    if (SandR)
      (posedge G *> (Q    +: D)) = (tplh$G$Q,    tphl$G$Q);
    if (SandRandCLK)
      ( D *> Q ) = (tplh$D$Q, tphl$D$Q );
    $setuphold(negedge G, posedge RN &&& (xSN == 1'b1), tsetup$RN$G,thold$RN$G, NOTIFIER);
    $width(negedge RN &&& (xSN == 1'b1), tminpwl$RN, 0, NOTIFIER);

    // timing checks 7
    $setuphold(negedge G &&& (SandR == 1), posedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $setuphold(negedge G &&& (SandR == 1), negedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $width(posedge G &&& (SandR == 1), tminpwh$G, 0, NOTIFIER);
    $period(posedge G &&& (SandR == 1), tperiod$G, NOTIFIER);
    if (D == 1'b0 && G == 1'b0 )
       (negedge  RN *> (Q +: 1'b1)) = ( tphl$RN$Q);
    if (D == 1'b1 && G == 1'b0 )
       (negedge  RN *> (Q +: 1'b1)) = ( tphl$RN$Q);
    if (D == 1'b1 && G == 1'b1 )
       (negedge  RN *> (Q +: 1'b1)) = (tplh$RN$Q, tphl$RN$Q);

   endspecify
endmodule //LATRQX3MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATRQX2MA10TR (Q, D, G, RN);
output  Q;
input  D, G, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

buf       XX0 (xRN, RN);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
not I3(clk,G);
buf I4(flgclk,G);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$Q   = 1.0,
      tphl$D$Q   = 1.0,
      tplh$G$Q   = 1.0,
      tphl$G$Q   = 1.0,
      tplh$RN$Q   = 1.0,
      tphl$RN$Q   = 1.0,
      tsetup$D$G = 1.0,
      thold$D$G  = 0.5,
      tsetup$D$RN = 1.0,
      thold$D$RN  = 0.5,
      tsetup$G$RN = 1.0,
      thold$G$RN  = 0.5,
      tsetup$RN$G = 1.0,
      thold$RN$G  = 0.5,
      tminpwl$RN    = 1.0,
      tminpwh$G  = 1.0,
      tperiod$G  = 1.0;
    // path delays
    if (SandR)
      (posedge G *> (Q    +: D)) = (tplh$G$Q,    tphl$G$Q);
    if (SandRandCLK)
      ( D *> Q ) = (tplh$D$Q, tphl$D$Q );
    $setuphold(negedge G, posedge RN &&& (xSN == 1'b1), tsetup$RN$G,thold$RN$G, NOTIFIER);
    $width(negedge RN &&& (xSN == 1'b1), tminpwl$RN, 0, NOTIFIER);

    // timing checks 7
    $setuphold(negedge G &&& (SandR == 1), posedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $setuphold(negedge G &&& (SandR == 1), negedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $width(posedge G &&& (SandR == 1), tminpwh$G, 0, NOTIFIER);
    $period(posedge G &&& (SandR == 1), tperiod$G, NOTIFIER);
    if (D == 1'b0 && G == 1'b0 )
       (negedge  RN *> (Q +: 1'b1)) = ( tphl$RN$Q);
    if (D == 1'b1 && G == 1'b0 )
       (negedge  RN *> (Q +: 1'b1)) = ( tphl$RN$Q);
    if (D == 1'b1 && G == 1'b1 )
       (negedge  RN *> (Q +: 1'b1)) = (tplh$RN$Q, tphl$RN$Q);

   endspecify
endmodule //LATRQX2MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATRQX1MA10TR (Q, D, G, RN);
output  Q;
input  D, G, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

buf       XX0 (xRN, RN);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
not I3(clk,G);
buf I4(flgclk,G);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$Q   = 1.0,
      tphl$D$Q   = 1.0,
      tplh$G$Q   = 1.0,
      tphl$G$Q   = 1.0,
      tplh$RN$Q   = 1.0,
      tphl$RN$Q   = 1.0,
      tsetup$D$G = 1.0,
      thold$D$G  = 0.5,
      tsetup$D$RN = 1.0,
      thold$D$RN  = 0.5,
      tsetup$G$RN = 1.0,
      thold$G$RN  = 0.5,
      tsetup$RN$G = 1.0,
      thold$RN$G  = 0.5,
      tminpwl$RN    = 1.0,
      tminpwh$G  = 1.0,
      tperiod$G  = 1.0;
    // path delays
    if (SandR)
      (posedge G *> (Q    +: D)) = (tplh$G$Q,    tphl$G$Q);
    if (SandRandCLK)
      ( D *> Q ) = (tplh$D$Q, tphl$D$Q );
    $setuphold(negedge G, posedge RN &&& (xSN == 1'b1), tsetup$RN$G,thold$RN$G, NOTIFIER);
    $width(negedge RN &&& (xSN == 1'b1), tminpwl$RN, 0, NOTIFIER);

    // timing checks 7
    $setuphold(negedge G &&& (SandR == 1), posedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $setuphold(negedge G &&& (SandR == 1), negedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $width(posedge G &&& (SandR == 1), tminpwh$G, 0, NOTIFIER);
    $period(posedge G &&& (SandR == 1), tperiod$G, NOTIFIER);
    if (D == 1'b0 && G == 1'b0 )
       (negedge  RN *> (Q +: 1'b1)) = ( tphl$RN$Q);
    if (D == 1'b1 && G == 1'b0 )
       (negedge  RN *> (Q +: 1'b1)) = ( tphl$RN$Q);
    if (D == 1'b1 && G == 1'b1 )
       (negedge  RN *> (Q +: 1'b1)) = (tplh$RN$Q, tphl$RN$Q);

   endspecify
endmodule //LATRQX1MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATRQX0P5MA10TR (Q, D, G, RN);
output  Q;
input  D, G, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

buf       XX0 (xRN, RN);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
not I3(clk,G);
buf I4(flgclk,G);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$Q   = 1.0,
      tphl$D$Q   = 1.0,
      tplh$G$Q   = 1.0,
      tphl$G$Q   = 1.0,
      tplh$RN$Q   = 1.0,
      tphl$RN$Q   = 1.0,
      tsetup$D$G = 1.0,
      thold$D$G  = 0.5,
      tsetup$D$RN = 1.0,
      thold$D$RN  = 0.5,
      tsetup$G$RN = 1.0,
      thold$G$RN  = 0.5,
      tsetup$RN$G = 1.0,
      thold$RN$G  = 0.5,
      tminpwl$RN    = 1.0,
      tminpwh$G  = 1.0,
      tperiod$G  = 1.0;
    // path delays
    if (SandR)
      (posedge G *> (Q    +: D)) = (tplh$G$Q,    tphl$G$Q);
    if (SandRandCLK)
      ( D *> Q ) = (tplh$D$Q, tphl$D$Q );
    $setuphold(negedge G, posedge RN &&& (xSN == 1'b1), tsetup$RN$G,thold$RN$G, NOTIFIER);
    $width(negedge RN &&& (xSN == 1'b1), tminpwl$RN, 0, NOTIFIER);

    // timing checks 7
    $setuphold(negedge G &&& (SandR == 1), posedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $setuphold(negedge G &&& (SandR == 1), negedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $width(posedge G &&& (SandR == 1), tminpwh$G, 0, NOTIFIER);
    $period(posedge G &&& (SandR == 1), tperiod$G, NOTIFIER);
    if (D == 1'b0 && G == 1'b0 )
       (negedge  RN *> (Q +: 1'b1)) = ( tphl$RN$Q);
    if (D == 1'b1 && G == 1'b0 )
       (negedge  RN *> (Q +: 1'b1)) = ( tphl$RN$Q);
    if (D == 1'b1 && G == 1'b1 )
       (negedge  RN *> (Q +: 1'b1)) = (tplh$RN$Q, tphl$RN$Q);

   endspecify
endmodule //LATRQX0P5MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATRPQNX4MA10TR (QN, D, G, R);
output  QN;
input  D, G, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

not       XX0 (xRN, R);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
not I3(clk,G);
buf I4(flgclk,G);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$QN   = 1.0,
      tphl$D$QN   = 1.0,
      tplh$G$QN   = 1.0,
      tphl$G$QN   = 1.0,
      tplh$R$QN   = 1.0,
      tphl$R$QN   = 1.0,
      tsetup$D$G = 1.0,
      thold$D$G  = 0.5,
      tsetup$D$R = 1.0,
      thold$D$R  = 0.5,
      tsetup$G$R = 1.0,
      thold$G$R  = 0.5,
      tsetup$R$G = 1.0,
      thold$R$G  = 0.5,
      tminpwh$R    = 1.0,
      tminpwh$G  = 1.0,
      tperiod$G  = 1.0;
    // path delays
    if (SandR)
      (posedge G *> (QN    -: D)) = (tplh$G$QN,    tphl$G$QN);
    if (SandRandCLK)
      ( D *> QN ) = (tplh$D$QN, tphl$D$QN );
    $setuphold(negedge G, negedge R, tsetup$R$G,thold$R$G, NOTIFIER);
    $width(posedge R, tminpwh$R, 0, NOTIFIER);
    // timing checks 2
    $setuphold(negedge G &&& (SandR == 1), posedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $setuphold(negedge G &&& (SandR == 1), negedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $width(posedge G &&& (SandR == 1), tminpwh$G, 0, NOTIFIER);
    $period(posedge G &&& (SandR == 1), tperiod$G, NOTIFIER);
    if (D == 1'b0 && G == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = ( tphl$R$QN);
    if (D == 1'b1 && G == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = ( tphl$R$QN);
    if (D == 1'b1 && G == 1'b1 )
       (posedge  R *> (QN -: 1'b1)) = (tplh$R$QN, tphl$R$QN);

   endspecify
endmodule //LATRPQNX4MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATRPQNX3MA10TR (QN, D, G, R);
output  QN;
input  D, G, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

not       XX0 (xRN, R);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
not I3(clk,G);
buf I4(flgclk,G);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$QN   = 1.0,
      tphl$D$QN   = 1.0,
      tplh$G$QN   = 1.0,
      tphl$G$QN   = 1.0,
      tplh$R$QN   = 1.0,
      tphl$R$QN   = 1.0,
      tsetup$D$G = 1.0,
      thold$D$G  = 0.5,
      tsetup$D$R = 1.0,
      thold$D$R  = 0.5,
      tsetup$G$R = 1.0,
      thold$G$R  = 0.5,
      tsetup$R$G = 1.0,
      thold$R$G  = 0.5,
      tminpwh$R    = 1.0,
      tminpwh$G  = 1.0,
      tperiod$G  = 1.0;
    // path delays
    if (SandR)
      (posedge G *> (QN    -: D)) = (tplh$G$QN,    tphl$G$QN);
    if (SandRandCLK)
      ( D *> QN ) = (tplh$D$QN, tphl$D$QN );
    $setuphold(negedge G, negedge R, tsetup$R$G,thold$R$G, NOTIFIER);
    $width(posedge R, tminpwh$R, 0, NOTIFIER);
    // timing checks 2
    $setuphold(negedge G &&& (SandR == 1), posedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $setuphold(negedge G &&& (SandR == 1), negedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $width(posedge G &&& (SandR == 1), tminpwh$G, 0, NOTIFIER);
    $period(posedge G &&& (SandR == 1), tperiod$G, NOTIFIER);
    if (D == 1'b0 && G == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = ( tphl$R$QN);
    if (D == 1'b1 && G == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = ( tphl$R$QN);
    if (D == 1'b1 && G == 1'b1 )
       (posedge  R *> (QN -: 1'b1)) = (tplh$R$QN, tphl$R$QN);

   endspecify
endmodule //LATRPQNX3MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATRPQNX2MA10TR (QN, D, G, R);
output  QN;
input  D, G, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

not       XX0 (xRN, R);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
not I3(clk,G);
buf I4(flgclk,G);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$QN   = 1.0,
      tphl$D$QN   = 1.0,
      tplh$G$QN   = 1.0,
      tphl$G$QN   = 1.0,
      tplh$R$QN   = 1.0,
      tphl$R$QN   = 1.0,
      tsetup$D$G = 1.0,
      thold$D$G  = 0.5,
      tsetup$D$R = 1.0,
      thold$D$R  = 0.5,
      tsetup$G$R = 1.0,
      thold$G$R  = 0.5,
      tsetup$R$G = 1.0,
      thold$R$G  = 0.5,
      tminpwh$R    = 1.0,
      tminpwh$G  = 1.0,
      tperiod$G  = 1.0;
    // path delays
    if (SandR)
      (posedge G *> (QN    -: D)) = (tplh$G$QN,    tphl$G$QN);
    if (SandRandCLK)
      ( D *> QN ) = (tplh$D$QN, tphl$D$QN );
    $setuphold(negedge G, negedge R, tsetup$R$G,thold$R$G, NOTIFIER);
    $width(posedge R, tminpwh$R, 0, NOTIFIER);
    // timing checks 2
    $setuphold(negedge G &&& (SandR == 1), posedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $setuphold(negedge G &&& (SandR == 1), negedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $width(posedge G &&& (SandR == 1), tminpwh$G, 0, NOTIFIER);
    $period(posedge G &&& (SandR == 1), tperiod$G, NOTIFIER);
    if (D == 1'b0 && G == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = ( tphl$R$QN);
    if (D == 1'b1 && G == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = ( tphl$R$QN);
    if (D == 1'b1 && G == 1'b1 )
       (posedge  R *> (QN -: 1'b1)) = (tplh$R$QN, tphl$R$QN);

   endspecify
endmodule //LATRPQNX2MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATRPQNX1MA10TR (QN, D, G, R);
output  QN;
input  D, G, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

not       XX0 (xRN, R);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
not I3(clk,G);
buf I4(flgclk,G);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$QN   = 1.0,
      tphl$D$QN   = 1.0,
      tplh$G$QN   = 1.0,
      tphl$G$QN   = 1.0,
      tplh$R$QN   = 1.0,
      tphl$R$QN   = 1.0,
      tsetup$D$G = 1.0,
      thold$D$G  = 0.5,
      tsetup$D$R = 1.0,
      thold$D$R  = 0.5,
      tsetup$G$R = 1.0,
      thold$G$R  = 0.5,
      tsetup$R$G = 1.0,
      thold$R$G  = 0.5,
      tminpwh$R    = 1.0,
      tminpwh$G  = 1.0,
      tperiod$G  = 1.0;
    // path delays
    if (SandR)
      (posedge G *> (QN    -: D)) = (tplh$G$QN,    tphl$G$QN);
    if (SandRandCLK)
      ( D *> QN ) = (tplh$D$QN, tphl$D$QN );
    $setuphold(negedge G, negedge R, tsetup$R$G,thold$R$G, NOTIFIER);
    $width(posedge R, tminpwh$R, 0, NOTIFIER);
    // timing checks 2
    $setuphold(negedge G &&& (SandR == 1), posedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $setuphold(negedge G &&& (SandR == 1), negedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $width(posedge G &&& (SandR == 1), tminpwh$G, 0, NOTIFIER);
    $period(posedge G &&& (SandR == 1), tperiod$G, NOTIFIER);
    if (D == 1'b0 && G == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = ( tphl$R$QN);
    if (D == 1'b1 && G == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = ( tphl$R$QN);
    if (D == 1'b1 && G == 1'b1 )
       (posedge  R *> (QN -: 1'b1)) = (tplh$R$QN, tphl$R$QN);

   endspecify
endmodule //LATRPQNX1MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATRPQNX0P5MA10TR (QN, D, G, R);
output  QN;
input  D, G, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

not       XX0 (xRN, R);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
not I3(clk,G);
buf I4(flgclk,G);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$QN   = 1.0,
      tphl$D$QN   = 1.0,
      tplh$G$QN   = 1.0,
      tphl$G$QN   = 1.0,
      tplh$R$QN   = 1.0,
      tphl$R$QN   = 1.0,
      tsetup$D$G = 1.0,
      thold$D$G  = 0.5,
      tsetup$D$R = 1.0,
      thold$D$R  = 0.5,
      tsetup$G$R = 1.0,
      thold$G$R  = 0.5,
      tsetup$R$G = 1.0,
      thold$R$G  = 0.5,
      tminpwh$R    = 1.0,
      tminpwh$G  = 1.0,
      tperiod$G  = 1.0;
    // path delays
    if (SandR)
      (posedge G *> (QN    -: D)) = (tplh$G$QN,    tphl$G$QN);
    if (SandRandCLK)
      ( D *> QN ) = (tplh$D$QN, tphl$D$QN );
    $setuphold(negedge G, negedge R, tsetup$R$G,thold$R$G, NOTIFIER);
    $width(posedge R, tminpwh$R, 0, NOTIFIER);
    // timing checks 2
    $setuphold(negedge G &&& (SandR == 1), posedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $setuphold(negedge G &&& (SandR == 1), negedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $width(posedge G &&& (SandR == 1), tminpwh$G, 0, NOTIFIER);
    $period(posedge G &&& (SandR == 1), tperiod$G, NOTIFIER);
    if (D == 1'b0 && G == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = ( tphl$R$QN);
    if (D == 1'b1 && G == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = ( tphl$R$QN);
    if (D == 1'b1 && G == 1'b1 )
       (posedge  R *> (QN -: 1'b1)) = (tplh$R$QN, tphl$R$QN);

   endspecify
endmodule //LATRPQNX0P5MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATQNX4MA10TR (QN, D, G);
output  QN;
input  D, G;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
not I3(clk,G);
buf I4(flgclk,G);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$QN   = 1.0,
      tphl$D$QN   = 1.0,
      tplh$G$QN   = 1.0,
      tphl$G$QN   = 1.0,
      tsetup$D$G = 1.0,
      thold$D$G  = 0.5,
      tminpwh$G  = 1.0,
      tperiod$G  = 1.0;
    // path delays
    if (SandR)
      (posedge G *> (QN    -: D)) = (tplh$G$QN,    tphl$G$QN);
    if (SandRandCLK)
      ( D *> QN ) = (tplh$D$QN, tphl$D$QN );
    // timing checks 2
    $setuphold(negedge G &&& (SandR == 1), posedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $setuphold(negedge G &&& (SandR == 1), negedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $width(posedge G &&& (SandR == 1), tminpwh$G, 0, NOTIFIER);
    $period(posedge G &&& (SandR == 1), tperiod$G, NOTIFIER);

   endspecify
endmodule //LATQNX4MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATQNX3MA10TR (QN, D, G);
output  QN;
input  D, G;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
not I3(clk,G);
buf I4(flgclk,G);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$QN   = 1.0,
      tphl$D$QN   = 1.0,
      tplh$G$QN   = 1.0,
      tphl$G$QN   = 1.0,
      tsetup$D$G = 1.0,
      thold$D$G  = 0.5,
      tminpwh$G  = 1.0,
      tperiod$G  = 1.0;
    // path delays
    if (SandR)
      (posedge G *> (QN    -: D)) = (tplh$G$QN,    tphl$G$QN);
    if (SandRandCLK)
      ( D *> QN ) = (tplh$D$QN, tphl$D$QN );
    // timing checks 2
    $setuphold(negedge G &&& (SandR == 1), posedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $setuphold(negedge G &&& (SandR == 1), negedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $width(posedge G &&& (SandR == 1), tminpwh$G, 0, NOTIFIER);
    $period(posedge G &&& (SandR == 1), tperiod$G, NOTIFIER);

   endspecify
endmodule //LATQNX3MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATQNX2MA10TR (QN, D, G);
output  QN;
input  D, G;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
not I3(clk,G);
buf I4(flgclk,G);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$QN   = 1.0,
      tphl$D$QN   = 1.0,
      tplh$G$QN   = 1.0,
      tphl$G$QN   = 1.0,
      tsetup$D$G = 1.0,
      thold$D$G  = 0.5,
      tminpwh$G  = 1.0,
      tperiod$G  = 1.0;
    // path delays
    if (SandR)
      (posedge G *> (QN    -: D)) = (tplh$G$QN,    tphl$G$QN);
    if (SandRandCLK)
      ( D *> QN ) = (tplh$D$QN, tphl$D$QN );
    // timing checks 2
    $setuphold(negedge G &&& (SandR == 1), posedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $setuphold(negedge G &&& (SandR == 1), negedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $width(posedge G &&& (SandR == 1), tminpwh$G, 0, NOTIFIER);
    $period(posedge G &&& (SandR == 1), tperiod$G, NOTIFIER);

   endspecify
endmodule //LATQNX2MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATQNX1MA10TR (QN, D, G);
output  QN;
input  D, G;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
not I3(clk,G);
buf I4(flgclk,G);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$QN   = 1.0,
      tphl$D$QN   = 1.0,
      tplh$G$QN   = 1.0,
      tphl$G$QN   = 1.0,
      tsetup$D$G = 1.0,
      thold$D$G  = 0.5,
      tminpwh$G  = 1.0,
      tperiod$G  = 1.0;
    // path delays
    if (SandR)
      (posedge G *> (QN    -: D)) = (tplh$G$QN,    tphl$G$QN);
    if (SandRandCLK)
      ( D *> QN ) = (tplh$D$QN, tphl$D$QN );
    // timing checks 2
    $setuphold(negedge G &&& (SandR == 1), posedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $setuphold(negedge G &&& (SandR == 1), negedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $width(posedge G &&& (SandR == 1), tminpwh$G, 0, NOTIFIER);
    $period(posedge G &&& (SandR == 1), tperiod$G, NOTIFIER);

   endspecify
endmodule //LATQNX1MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATQNX0P5MA10TR (QN, D, G);
output  QN;
input  D, G;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
not I3(clk,G);
buf I4(flgclk,G);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$QN   = 1.0,
      tphl$D$QN   = 1.0,
      tplh$G$QN   = 1.0,
      tphl$G$QN   = 1.0,
      tsetup$D$G = 1.0,
      thold$D$G  = 0.5,
      tminpwh$G  = 1.0,
      tperiod$G  = 1.0;
    // path delays
    if (SandR)
      (posedge G *> (QN    -: D)) = (tplh$G$QN,    tphl$G$QN);
    if (SandRandCLK)
      ( D *> QN ) = (tplh$D$QN, tphl$D$QN );
    // timing checks 2
    $setuphold(negedge G &&& (SandR == 1), posedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $setuphold(negedge G &&& (SandR == 1), negedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $width(posedge G &&& (SandR == 1), tminpwh$G, 0, NOTIFIER);
    $period(posedge G &&& (SandR == 1), tperiod$G, NOTIFIER);

   endspecify
endmodule //LATQNX0P5MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATQX3MA10TR (Q, D, G);
output  Q;
input  D, G;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
not I3(clk,G);
buf I4(flgclk,G);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$Q   = 1.0,
      tphl$D$Q   = 1.0,
      tplh$G$Q   = 1.0,
      tphl$G$Q   = 1.0,
      tsetup$D$G = 1.0,
      thold$D$G  = 0.5,
      tminpwh$G  = 1.0,
      tperiod$G  = 1.0;
    // path delays
    if (SandR)
      (posedge G *> (Q    +: D)) = (tplh$G$Q,    tphl$G$Q);
    if (SandRandCLK)
      ( D *> Q ) = (tplh$D$Q, tphl$D$Q );

    // timing checks 7
    $setuphold(negedge G &&& (SandR == 1), posedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $setuphold(negedge G &&& (SandR == 1), negedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $width(posedge G &&& (SandR == 1), tminpwh$G, 0, NOTIFIER);
    $period(posedge G &&& (SandR == 1), tperiod$G, NOTIFIER);

   endspecify
endmodule //LATQX3MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATQX2MA10TR (Q, D, G);
output  Q;
input  D, G;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
not I3(clk,G);
buf I4(flgclk,G);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$Q   = 1.0,
      tphl$D$Q   = 1.0,
      tplh$G$Q   = 1.0,
      tphl$G$Q   = 1.0,
      tsetup$D$G = 1.0,
      thold$D$G  = 0.5,
      tminpwh$G  = 1.0,
      tperiod$G  = 1.0;
    // path delays
    if (SandR)
      (posedge G *> (Q    +: D)) = (tplh$G$Q,    tphl$G$Q);
    if (SandRandCLK)
      ( D *> Q ) = (tplh$D$Q, tphl$D$Q );

    // timing checks 7
    $setuphold(negedge G &&& (SandR == 1), posedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $setuphold(negedge G &&& (SandR == 1), negedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $width(posedge G &&& (SandR == 1), tminpwh$G, 0, NOTIFIER);
    $period(posedge G &&& (SandR == 1), tperiod$G, NOTIFIER);

   endspecify
endmodule //LATQX2MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATQX1MA10TR (Q, D, G);
output  Q;
input  D, G;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
not I3(clk,G);
buf I4(flgclk,G);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$Q   = 1.0,
      tphl$D$Q   = 1.0,
      tplh$G$Q   = 1.0,
      tphl$G$Q   = 1.0,
      tsetup$D$G = 1.0,
      thold$D$G  = 0.5,
      tminpwh$G  = 1.0,
      tperiod$G  = 1.0;
    // path delays
    if (SandR)
      (posedge G *> (Q    +: D)) = (tplh$G$Q,    tphl$G$Q);
    if (SandRandCLK)
      ( D *> Q ) = (tplh$D$Q, tphl$D$Q );

    // timing checks 7
    $setuphold(negedge G &&& (SandR == 1), posedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $setuphold(negedge G &&& (SandR == 1), negedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $width(posedge G &&& (SandR == 1), tminpwh$G, 0, NOTIFIER);
    $period(posedge G &&& (SandR == 1), tperiod$G, NOTIFIER);

   endspecify
endmodule //LATQX1MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATQX0P5MA10TR (Q, D, G);
output  Q;
input  D, G;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
not I3(clk,G);
buf I4(flgclk,G);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$Q   = 1.0,
      tphl$D$Q   = 1.0,
      tplh$G$Q   = 1.0,
      tphl$G$Q   = 1.0,
      tsetup$D$G = 1.0,
      thold$D$G  = 0.5,
      tminpwh$G  = 1.0,
      tperiod$G  = 1.0;
    // path delays
    if (SandR)
      (posedge G *> (Q    +: D)) = (tplh$G$Q,    tphl$G$Q);
    if (SandRandCLK)
      ( D *> Q ) = (tplh$D$Q, tphl$D$Q );

    // timing checks 7
    $setuphold(negedge G &&& (SandR == 1), posedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $setuphold(negedge G &&& (SandR == 1), negedge D, tsetup$D$G,thold$D$G, NOTIFIER);
    $width(posedge G &&& (SandR == 1), tminpwh$G, 0, NOTIFIER);
    $period(posedge G &&& (SandR == 1), tperiod$G, NOTIFIER);

   endspecify
endmodule //LATQX0P5MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATNSQNX4MA10TR (QN, D, GN, SN);
output  QN;
input  D, GN, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

buf       XX0 (xSN, SN);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$QN   = 1.0,
      tphl$D$QN   = 1.0,
      tplh$GN$QN   = 1.0,
      tphl$GN$QN   = 1.0,
      tplh$SN$QN   = 1.0,
      tphl$SN$QN   = 1.0,
      tsetup$D$GN = 1.0,
      thold$D$GN  = 0.5,
      tsetup$D$SN = 1.0,
      thold$D$SN  = 0.5,
      tsetup$GN$SN = 1.0,
      thold$GN$SN  = 0.5,
      tsetup$SN$GN = 1.0,
      thold$SN$GN  = 0.5,
      tminpwl$SN  = 1.0,
      tminpwl$GN  = 1.0,
      tperiod$GN  = 1.0;
    // path delays
    if (SandR)
      (negedge GN *> (QN    -: D)) = (tplh$GN$QN,    tphl$GN$QN);
    if (SandRandCLK)
      ( D *> QN ) = (tplh$D$QN, tphl$D$QN );
    $setuphold(posedge GN, posedge SN, tsetup$SN$GN,thold$SN$GN, NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    // timing checks 1
    $setuphold(posedge GN &&& (SandR == 1), posedge D, tsetup$D$GN,thold$D$GN, NOTIFIER);
    $setuphold(posedge GN &&& (SandR == 1), negedge D, tsetup$D$GN,thold$D$GN, NOTIFIER);
    $width(negedge GN &&& (SandR == 1), tminpwl$GN, 0, NOTIFIER);
    $period(posedge GN &&& (SandR == 1), tperiod$GN, NOTIFIER);
    if (D == 1'b0 && GN == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN);
    if (D == 1'b0 && GN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN);
    if (D == 1'b1 && GN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN);

   endspecify
endmodule //LATNSQNX4MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATNSQNX3MA10TR (QN, D, GN, SN);
output  QN;
input  D, GN, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

buf       XX0 (xSN, SN);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$QN   = 1.0,
      tphl$D$QN   = 1.0,
      tplh$GN$QN   = 1.0,
      tphl$GN$QN   = 1.0,
      tplh$SN$QN   = 1.0,
      tphl$SN$QN   = 1.0,
      tsetup$D$GN = 1.0,
      thold$D$GN  = 0.5,
      tsetup$D$SN = 1.0,
      thold$D$SN  = 0.5,
      tsetup$GN$SN = 1.0,
      thold$GN$SN  = 0.5,
      tsetup$SN$GN = 1.0,
      thold$SN$GN  = 0.5,
      tminpwl$SN  = 1.0,
      tminpwl$GN  = 1.0,
      tperiod$GN  = 1.0;
    // path delays
    if (SandR)
      (negedge GN *> (QN    -: D)) = (tplh$GN$QN,    tphl$GN$QN);
    if (SandRandCLK)
      ( D *> QN ) = (tplh$D$QN, tphl$D$QN );
    $setuphold(posedge GN, posedge SN, tsetup$SN$GN,thold$SN$GN, NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    // timing checks 1
    $setuphold(posedge GN &&& (SandR == 1), posedge D, tsetup$D$GN,thold$D$GN, NOTIFIER);
    $setuphold(posedge GN &&& (SandR == 1), negedge D, tsetup$D$GN,thold$D$GN, NOTIFIER);
    $width(negedge GN &&& (SandR == 1), tminpwl$GN, 0, NOTIFIER);
    $period(posedge GN &&& (SandR == 1), tperiod$GN, NOTIFIER);
    if (D == 1'b0 && GN == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN);
    if (D == 1'b0 && GN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN);
    if (D == 1'b1 && GN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN);

   endspecify
endmodule //LATNSQNX3MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATNSQNX2MA10TR (QN, D, GN, SN);
output  QN;
input  D, GN, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

buf       XX0 (xSN, SN);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$QN   = 1.0,
      tphl$D$QN   = 1.0,
      tplh$GN$QN   = 1.0,
      tphl$GN$QN   = 1.0,
      tplh$SN$QN   = 1.0,
      tphl$SN$QN   = 1.0,
      tsetup$D$GN = 1.0,
      thold$D$GN  = 0.5,
      tsetup$D$SN = 1.0,
      thold$D$SN  = 0.5,
      tsetup$GN$SN = 1.0,
      thold$GN$SN  = 0.5,
      tsetup$SN$GN = 1.0,
      thold$SN$GN  = 0.5,
      tminpwl$SN  = 1.0,
      tminpwl$GN  = 1.0,
      tperiod$GN  = 1.0;
    // path delays
    if (SandR)
      (negedge GN *> (QN    -: D)) = (tplh$GN$QN,    tphl$GN$QN);
    if (SandRandCLK)
      ( D *> QN ) = (tplh$D$QN, tphl$D$QN );
    $setuphold(posedge GN, posedge SN, tsetup$SN$GN,thold$SN$GN, NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    // timing checks 1
    $setuphold(posedge GN &&& (SandR == 1), posedge D, tsetup$D$GN,thold$D$GN, NOTIFIER);
    $setuphold(posedge GN &&& (SandR == 1), negedge D, tsetup$D$GN,thold$D$GN, NOTIFIER);
    $width(negedge GN &&& (SandR == 1), tminpwl$GN, 0, NOTIFIER);
    $period(posedge GN &&& (SandR == 1), tperiod$GN, NOTIFIER);
    if (D == 1'b0 && GN == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN);
    if (D == 1'b0 && GN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN);
    if (D == 1'b1 && GN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN);

   endspecify
endmodule //LATNSQNX2MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATNSQNX1MA10TR (QN, D, GN, SN);
output  QN;
input  D, GN, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

buf       XX0 (xSN, SN);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$QN   = 1.0,
      tphl$D$QN   = 1.0,
      tplh$GN$QN   = 1.0,
      tphl$GN$QN   = 1.0,
      tplh$SN$QN   = 1.0,
      tphl$SN$QN   = 1.0,
      tsetup$D$GN = 1.0,
      thold$D$GN  = 0.5,
      tsetup$D$SN = 1.0,
      thold$D$SN  = 0.5,
      tsetup$GN$SN = 1.0,
      thold$GN$SN  = 0.5,
      tsetup$SN$GN = 1.0,
      thold$SN$GN  = 0.5,
      tminpwl$SN  = 1.0,
      tminpwl$GN  = 1.0,
      tperiod$GN  = 1.0;
    // path delays
    if (SandR)
      (negedge GN *> (QN    -: D)) = (tplh$GN$QN,    tphl$GN$QN);
    if (SandRandCLK)
      ( D *> QN ) = (tplh$D$QN, tphl$D$QN );
    $setuphold(posedge GN, posedge SN, tsetup$SN$GN,thold$SN$GN, NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    // timing checks 1
    $setuphold(posedge GN &&& (SandR == 1), posedge D, tsetup$D$GN,thold$D$GN, NOTIFIER);
    $setuphold(posedge GN &&& (SandR == 1), negedge D, tsetup$D$GN,thold$D$GN, NOTIFIER);
    $width(negedge GN &&& (SandR == 1), tminpwl$GN, 0, NOTIFIER);
    $period(posedge GN &&& (SandR == 1), tperiod$GN, NOTIFIER);
    if (D == 1'b0 && GN == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN);
    if (D == 1'b0 && GN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN);
    if (D == 1'b1 && GN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN);

   endspecify
endmodule //LATNSQNX1MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATNSQNX0P5MA10TR (QN, D, GN, SN);
output  QN;
input  D, GN, SN;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

buf       XX0 (xSN, SN);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$QN   = 1.0,
      tphl$D$QN   = 1.0,
      tplh$GN$QN   = 1.0,
      tphl$GN$QN   = 1.0,
      tplh$SN$QN   = 1.0,
      tphl$SN$QN   = 1.0,
      tsetup$D$GN = 1.0,
      thold$D$GN  = 0.5,
      tsetup$D$SN = 1.0,
      thold$D$SN  = 0.5,
      tsetup$GN$SN = 1.0,
      thold$GN$SN  = 0.5,
      tsetup$SN$GN = 1.0,
      thold$SN$GN  = 0.5,
      tminpwl$SN  = 1.0,
      tminpwl$GN  = 1.0,
      tperiod$GN  = 1.0;
    // path delays
    if (SandR)
      (negedge GN *> (QN    -: D)) = (tplh$GN$QN,    tphl$GN$QN);
    if (SandRandCLK)
      ( D *> QN ) = (tplh$D$QN, tphl$D$QN );
    $setuphold(posedge GN, posedge SN, tsetup$SN$GN,thold$SN$GN, NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    // timing checks 1
    $setuphold(posedge GN &&& (SandR == 1), posedge D, tsetup$D$GN,thold$D$GN, NOTIFIER);
    $setuphold(posedge GN &&& (SandR == 1), negedge D, tsetup$D$GN,thold$D$GN, NOTIFIER);
    $width(negedge GN &&& (SandR == 1), tminpwl$GN, 0, NOTIFIER);
    $period(posedge GN &&& (SandR == 1), tperiod$GN, NOTIFIER);
    if (D == 1'b0 && GN == 1'b0 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN, tphl$SN$QN);
    if (D == 1'b0 && GN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN);
    if (D == 1'b1 && GN == 1'b1 )
       (negedge  SN *> (QN -: 1'b1)) = (tplh$SN$QN);

   endspecify
endmodule //LATNSQNX0P5MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATNSPQX3MA10TR (Q, D, GN, S);
output  Q;
input  D, GN, S;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

not       XX0 (xSN, S);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$Q   = 1.0,
      tphl$D$Q   = 1.0,
      tplh$GN$Q   = 1.0,
      tphl$GN$Q   = 1.0,
      tplh$S$Q   = 1.0,
      tphl$S$Q   = 1.0,
      tsetup$D$GN = 1.0,
      thold$D$GN  = 0.5,
      tsetup$D$S = 1.0,
      thold$D$S  = 0.5,
      tsetup$GN$S = 1.0,
      thold$GN$S  = 0.5,
      tsetup$S$GN = 1.0,
      thold$S$GN  = 0.5,
      tminpwh$S    = 1.0,
      tminpwl$GN  = 1.0,
      tperiod$GN  = 1.0;
    // path delays
    if (SandR)
      (negedge GN *> (Q    +: D)) = (tplh$GN$Q,    tphl$GN$Q);
    if (SandRandCLK)
      ( D *> Q ) = (tplh$D$Q, tphl$D$Q );

    // timing checks 4
    $setuphold(posedge GN &&& (SandR == 1), posedge D, tsetup$D$GN,thold$D$GN, NOTIFIER);
    $setuphold(posedge GN &&& (SandR == 1), negedge D, tsetup$D$GN,thold$D$GN, NOTIFIER); 
    $setuphold(posedge GN, negedge S, tsetup$S$GN, thold$S$GN, NOTIFIER);
    $width(posedge S, tminpwh$S, 0, NOTIFIER);
    $width(negedge GN &&& (SandR == 1), tminpwl$GN, 0, NOTIFIER);
    $period(negedge GN &&& (SandR == 1), tperiod$GN, NOTIFIER);

    if (D == 1'b0 && GN == 1'b0 )
       (posedge  S *> (Q +: 1'b1)) = (tplh$S$Q, tphl$S$Q);
    if (D == 1'b0 && GN == 1'b1 )
       (posedge  S *> (Q +: 1'b1)) = ( tphl$S$Q);
    if (D == 1'b1 && GN == 1'b1 )
       (posedge  S *> (Q +: 1'b1)) = ( tphl$S$Q);

   endspecify
endmodule //LATNSPQX3MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATNSPQX2MA10TR (Q, D, GN, S);
output  Q;
input  D, GN, S;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

not       XX0 (xSN, S);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$Q   = 1.0,
      tphl$D$Q   = 1.0,
      tplh$GN$Q   = 1.0,
      tphl$GN$Q   = 1.0,
      tplh$S$Q   = 1.0,
      tphl$S$Q   = 1.0,
      tsetup$D$GN = 1.0,
      thold$D$GN  = 0.5,
      tsetup$D$S = 1.0,
      thold$D$S  = 0.5,
      tsetup$GN$S = 1.0,
      thold$GN$S  = 0.5,
      tsetup$S$GN = 1.0,
      thold$S$GN  = 0.5,
      tminpwh$S    = 1.0,
      tminpwl$GN  = 1.0,
      tperiod$GN  = 1.0;
    // path delays
    if (SandR)
      (negedge GN *> (Q    +: D)) = (tplh$GN$Q,    tphl$GN$Q);
    if (SandRandCLK)
      ( D *> Q ) = (tplh$D$Q, tphl$D$Q );

    // timing checks 4
    $setuphold(posedge GN &&& (SandR == 1), posedge D, tsetup$D$GN,thold$D$GN, NOTIFIER);
    $setuphold(posedge GN &&& (SandR == 1), negedge D, tsetup$D$GN,thold$D$GN, NOTIFIER); 
    $setuphold(posedge GN, negedge S, tsetup$S$GN, thold$S$GN, NOTIFIER);
    $width(posedge S, tminpwh$S, 0, NOTIFIER);
    $width(negedge GN &&& (SandR == 1), tminpwl$GN, 0, NOTIFIER);
    $period(negedge GN &&& (SandR == 1), tperiod$GN, NOTIFIER);

    if (D == 1'b0 && GN == 1'b0 )
       (posedge  S *> (Q +: 1'b1)) = (tplh$S$Q, tphl$S$Q);
    if (D == 1'b0 && GN == 1'b1 )
       (posedge  S *> (Q +: 1'b1)) = ( tphl$S$Q);
    if (D == 1'b1 && GN == 1'b1 )
       (posedge  S *> (Q +: 1'b1)) = ( tphl$S$Q);

   endspecify
endmodule //LATNSPQX2MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATNSPQX1MA10TR (Q, D, GN, S);
output  Q;
input  D, GN, S;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

not       XX0 (xSN, S);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$Q   = 1.0,
      tphl$D$Q   = 1.0,
      tplh$GN$Q   = 1.0,
      tphl$GN$Q   = 1.0,
      tplh$S$Q   = 1.0,
      tphl$S$Q   = 1.0,
      tsetup$D$GN = 1.0,
      thold$D$GN  = 0.5,
      tsetup$D$S = 1.0,
      thold$D$S  = 0.5,
      tsetup$GN$S = 1.0,
      thold$GN$S  = 0.5,
      tsetup$S$GN = 1.0,
      thold$S$GN  = 0.5,
      tminpwh$S    = 1.0,
      tminpwl$GN  = 1.0,
      tperiod$GN  = 1.0;
    // path delays
    if (SandR)
      (negedge GN *> (Q    +: D)) = (tplh$GN$Q,    tphl$GN$Q);
    if (SandRandCLK)
      ( D *> Q ) = (tplh$D$Q, tphl$D$Q );

    // timing checks 4
    $setuphold(posedge GN &&& (SandR == 1), posedge D, tsetup$D$GN,thold$D$GN, NOTIFIER);
    $setuphold(posedge GN &&& (SandR == 1), negedge D, tsetup$D$GN,thold$D$GN, NOTIFIER); 
    $setuphold(posedge GN, negedge S, tsetup$S$GN, thold$S$GN, NOTIFIER);
    $width(posedge S, tminpwh$S, 0, NOTIFIER);
    $width(negedge GN &&& (SandR == 1), tminpwl$GN, 0, NOTIFIER);
    $period(negedge GN &&& (SandR == 1), tperiod$GN, NOTIFIER);

    if (D == 1'b0 && GN == 1'b0 )
       (posedge  S *> (Q +: 1'b1)) = (tplh$S$Q, tphl$S$Q);
    if (D == 1'b0 && GN == 1'b1 )
       (posedge  S *> (Q +: 1'b1)) = ( tphl$S$Q);
    if (D == 1'b1 && GN == 1'b1 )
       (posedge  S *> (Q +: 1'b1)) = ( tphl$S$Q);

   endspecify
endmodule //LATNSPQX1MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATNSPQX0P5MA10TR (Q, D, GN, S);
output  Q;
input  D, GN, S;
reg NOTIFIER;
supply1 xRN;
supply1 dRN;

not       XX0 (xSN, S);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$Q   = 1.0,
      tphl$D$Q   = 1.0,
      tplh$GN$Q   = 1.0,
      tphl$GN$Q   = 1.0,
      tplh$S$Q   = 1.0,
      tphl$S$Q   = 1.0,
      tsetup$D$GN = 1.0,
      thold$D$GN  = 0.5,
      tsetup$D$S = 1.0,
      thold$D$S  = 0.5,
      tsetup$GN$S = 1.0,
      thold$GN$S  = 0.5,
      tsetup$S$GN = 1.0,
      thold$S$GN  = 0.5,
      tminpwh$S    = 1.0,
      tminpwl$GN  = 1.0,
      tperiod$GN  = 1.0;
    // path delays
    if (SandR)
      (negedge GN *> (Q    +: D)) = (tplh$GN$Q,    tphl$GN$Q);
    if (SandRandCLK)
      ( D *> Q ) = (tplh$D$Q, tphl$D$Q );

    // timing checks 4
    $setuphold(posedge GN &&& (SandR == 1), posedge D, tsetup$D$GN,thold$D$GN, NOTIFIER);
    $setuphold(posedge GN &&& (SandR == 1), negedge D, tsetup$D$GN,thold$D$GN, NOTIFIER); 
    $setuphold(posedge GN, negedge S, tsetup$S$GN, thold$S$GN, NOTIFIER);
    $width(posedge S, tminpwh$S, 0, NOTIFIER);
    $width(negedge GN &&& (SandR == 1), tminpwl$GN, 0, NOTIFIER);
    $period(negedge GN &&& (SandR == 1), tperiod$GN, NOTIFIER);

    if (D == 1'b0 && GN == 1'b0 )
       (posedge  S *> (Q +: 1'b1)) = (tplh$S$Q, tphl$S$Q);
    if (D == 1'b0 && GN == 1'b1 )
       (posedge  S *> (Q +: 1'b1)) = ( tphl$S$Q);
    if (D == 1'b1 && GN == 1'b1 )
       (posedge  S *> (Q +: 1'b1)) = ( tphl$S$Q);

   endspecify
endmodule //LATNSPQX0P5MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATNRQX3MA10TR (Q, D, GN, RN);
output  Q;
input  D, GN, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

buf       XX0 (xRN, RN);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$Q   = 1.0,
      tphl$D$Q   = 1.0,
      tplh$GN$Q   = 1.0,
      tphl$GN$Q   = 1.0,
      tplh$RN$Q   = 1.0,
      tphl$RN$Q   = 1.0,
      tsetup$D$GN = 1.0,
      thold$D$GN  = 0.5,
      tsetup$D$RN = 1.0,
      thold$D$RN  = 0.5,
      tsetup$GN$RN = 1.0,
      thold$GN$RN  = 0.5,
      tsetup$RN$GN = 1.0,
      thold$RN$GN  = 0.5,
      tminpwl$RN    = 1.0,
      tminpwl$GN  = 1.0,
      tperiod$GN  = 1.0;
    // path delays
    if (SandR)
      (negedge GN *> (Q    +: D)) = (tplh$GN$Q,    tphl$GN$Q);
    if (SandRandCLK)
      ( D *> Q ) = (tplh$D$Q, tphl$D$Q );
    $setuphold(posedge GN, posedge RN &&& (xSN == 1'b1), tsetup$RN$GN,thold$RN$GN, NOTIFIER);
    $width(negedge RN &&& (xSN == 1'b1), tminpwl$RN, 0, NOTIFIER);

    // timing checks 4
    $setuphold(posedge GN &&& (SandR == 1), posedge D, tsetup$D$GN,thold$D$GN, NOTIFIER);
    $setuphold(posedge GN &&& (SandR == 1), negedge D, tsetup$D$GN,thold$D$GN, NOTIFIER); 
    $width(negedge GN &&& (SandR == 1), tminpwl$GN, 0, NOTIFIER);
    $period(negedge GN &&& (SandR == 1), tperiod$GN, NOTIFIER);

    if (D == 1'b0 && GN == 1'b1 )
       (negedge  RN *> (Q +: 1'b1)) = (tplh$RN$Q);
    if (D == 1'b1 && GN == 1'b0 )
       (negedge  RN *> (Q +: 1'b1)) = (tplh$RN$Q, tphl$RN$Q);
    if (D == 1'b1 && GN == 1'b1 )
       (negedge  RN *> (Q +: 1'b1)) = (tplh$RN$Q);

   endspecify
endmodule //LATNRQX3MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATNRQX2MA10TR (Q, D, GN, RN);
output  Q;
input  D, GN, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

buf       XX0 (xRN, RN);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$Q   = 1.0,
      tphl$D$Q   = 1.0,
      tplh$GN$Q   = 1.0,
      tphl$GN$Q   = 1.0,
      tplh$RN$Q   = 1.0,
      tphl$RN$Q   = 1.0,
      tsetup$D$GN = 1.0,
      thold$D$GN  = 0.5,
      tsetup$D$RN = 1.0,
      thold$D$RN  = 0.5,
      tsetup$GN$RN = 1.0,
      thold$GN$RN  = 0.5,
      tsetup$RN$GN = 1.0,
      thold$RN$GN  = 0.5,
      tminpwl$RN    = 1.0,
      tminpwl$GN  = 1.0,
      tperiod$GN  = 1.0;
    // path delays
    if (SandR)
      (negedge GN *> (Q    +: D)) = (tplh$GN$Q,    tphl$GN$Q);
    if (SandRandCLK)
      ( D *> Q ) = (tplh$D$Q, tphl$D$Q );
    $setuphold(posedge GN, posedge RN &&& (xSN == 1'b1), tsetup$RN$GN,thold$RN$GN, NOTIFIER);
    $width(negedge RN &&& (xSN == 1'b1), tminpwl$RN, 0, NOTIFIER);

    // timing checks 4
    $setuphold(posedge GN &&& (SandR == 1), posedge D, tsetup$D$GN,thold$D$GN, NOTIFIER);
    $setuphold(posedge GN &&& (SandR == 1), negedge D, tsetup$D$GN,thold$D$GN, NOTIFIER); 
    $width(negedge GN &&& (SandR == 1), tminpwl$GN, 0, NOTIFIER);
    $period(negedge GN &&& (SandR == 1), tperiod$GN, NOTIFIER);

    if (D == 1'b0 && GN == 1'b1 )
       (negedge  RN *> (Q +: 1'b1)) = (tplh$RN$Q);
    if (D == 1'b1 && GN == 1'b0 )
       (negedge  RN *> (Q +: 1'b1)) = (tplh$RN$Q, tphl$RN$Q);
    if (D == 1'b1 && GN == 1'b1 )
       (negedge  RN *> (Q +: 1'b1)) = (tplh$RN$Q);

   endspecify
endmodule //LATNRQX2MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATNRQX1MA10TR (Q, D, GN, RN);
output  Q;
input  D, GN, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

buf       XX0 (xRN, RN);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$Q   = 1.0,
      tphl$D$Q   = 1.0,
      tplh$GN$Q   = 1.0,
      tphl$GN$Q   = 1.0,
      tplh$RN$Q   = 1.0,
      tphl$RN$Q   = 1.0,
      tsetup$D$GN = 1.0,
      thold$D$GN  = 0.5,
      tsetup$D$RN = 1.0,
      thold$D$RN  = 0.5,
      tsetup$GN$RN = 1.0,
      thold$GN$RN  = 0.5,
      tsetup$RN$GN = 1.0,
      thold$RN$GN  = 0.5,
      tminpwl$RN    = 1.0,
      tminpwl$GN  = 1.0,
      tperiod$GN  = 1.0;
    // path delays
    if (SandR)
      (negedge GN *> (Q    +: D)) = (tplh$GN$Q,    tphl$GN$Q);
    if (SandRandCLK)
      ( D *> Q ) = (tplh$D$Q, tphl$D$Q );
    $setuphold(posedge GN, posedge RN &&& (xSN == 1'b1), tsetup$RN$GN,thold$RN$GN, NOTIFIER);
    $width(negedge RN &&& (xSN == 1'b1), tminpwl$RN, 0, NOTIFIER);

    // timing checks 4
    $setuphold(posedge GN &&& (SandR == 1), posedge D, tsetup$D$GN,thold$D$GN, NOTIFIER);
    $setuphold(posedge GN &&& (SandR == 1), negedge D, tsetup$D$GN,thold$D$GN, NOTIFIER); 
    $width(negedge GN &&& (SandR == 1), tminpwl$GN, 0, NOTIFIER);
    $period(negedge GN &&& (SandR == 1), tperiod$GN, NOTIFIER);

    if (D == 1'b0 && GN == 1'b1 )
       (negedge  RN *> (Q +: 1'b1)) = (tplh$RN$Q);
    if (D == 1'b1 && GN == 1'b0 )
       (negedge  RN *> (Q +: 1'b1)) = (tplh$RN$Q, tphl$RN$Q);
    if (D == 1'b1 && GN == 1'b1 )
       (negedge  RN *> (Q +: 1'b1)) = (tplh$RN$Q);

   endspecify
endmodule //LATNRQX1MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATNRQX0P5MA10TR (Q, D, GN, RN);
output  Q;
input  D, GN, RN;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

buf       XX0 (xRN, RN);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$Q   = 1.0,
      tphl$D$Q   = 1.0,
      tplh$GN$Q   = 1.0,
      tphl$GN$Q   = 1.0,
      tplh$RN$Q   = 1.0,
      tphl$RN$Q   = 1.0,
      tsetup$D$GN = 1.0,
      thold$D$GN  = 0.5,
      tsetup$D$RN = 1.0,
      thold$D$RN  = 0.5,
      tsetup$GN$RN = 1.0,
      thold$GN$RN  = 0.5,
      tsetup$RN$GN = 1.0,
      thold$RN$GN  = 0.5,
      tminpwl$RN    = 1.0,
      tminpwl$GN  = 1.0,
      tperiod$GN  = 1.0;
    // path delays
    if (SandR)
      (negedge GN *> (Q    +: D)) = (tplh$GN$Q,    tphl$GN$Q);
    if (SandRandCLK)
      ( D *> Q ) = (tplh$D$Q, tphl$D$Q );
    $setuphold(posedge GN, posedge RN &&& (xSN == 1'b1), tsetup$RN$GN,thold$RN$GN, NOTIFIER);
    $width(negedge RN &&& (xSN == 1'b1), tminpwl$RN, 0, NOTIFIER);

    // timing checks 4
    $setuphold(posedge GN &&& (SandR == 1), posedge D, tsetup$D$GN,thold$D$GN, NOTIFIER);
    $setuphold(posedge GN &&& (SandR == 1), negedge D, tsetup$D$GN,thold$D$GN, NOTIFIER); 
    $width(negedge GN &&& (SandR == 1), tminpwl$GN, 0, NOTIFIER);
    $period(negedge GN &&& (SandR == 1), tperiod$GN, NOTIFIER);

    if (D == 1'b0 && GN == 1'b1 )
       (negedge  RN *> (Q +: 1'b1)) = (tplh$RN$Q);
    if (D == 1'b1 && GN == 1'b0 )
       (negedge  RN *> (Q +: 1'b1)) = (tplh$RN$Q, tphl$RN$Q);
    if (D == 1'b1 && GN == 1'b1 )
       (negedge  RN *> (Q +: 1'b1)) = (tplh$RN$Q);

   endspecify
endmodule //LATNRQX0P5MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATNRPQNX4MA10TR (QN, D, GN, R);
output  QN;
input  D, GN, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

not       XX0 (xRN, R);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$QN   = 1.0,
      tphl$D$QN   = 1.0,
      tplh$GN$QN   = 1.0,
      tphl$GN$QN   = 1.0,
      tplh$R$QN   = 1.0,
      tphl$R$QN   = 1.0,
      tsetup$D$GN = 1.0,
      thold$D$GN  = 0.5,
      tsetup$D$R = 1.0,
      thold$D$R  = 0.5,
      tsetup$GN$R = 1.0,
      thold$GN$R  = 0.5,
      tsetup$R$GN = 1.0,
      thold$R$GN  = 0.5,
      tminpwh$R    = 1.0,
      tminpwl$GN  = 1.0,
      tperiod$GN  = 1.0;
    // path delays
    if (SandR)
      (negedge GN *> (QN    -: D)) = (tplh$GN$QN,    tphl$GN$QN);
    if (SandRandCLK)
      ( D *> QN ) = (tplh$D$QN, tphl$D$QN );
    $setuphold(posedge GN, negedge R, tsetup$R$GN,thold$R$GN, NOTIFIER);
    $width(posedge R, tminpwh$R, 0, NOTIFIER);
    // timing checks 1
    $setuphold(posedge GN &&& (SandR == 1), posedge D, tsetup$D$GN,thold$D$GN, NOTIFIER);
    $setuphold(posedge GN &&& (SandR == 1), negedge D, tsetup$D$GN,thold$D$GN, NOTIFIER);
    $width(negedge GN &&& (SandR == 1), tminpwl$GN, 0, NOTIFIER);
    $period(posedge GN &&& (SandR == 1), tperiod$GN, NOTIFIER);
    if (D == 1'b0 && GN == 1'b1 )
       (posedge  R *> (QN -: 1'b0)) = ( tphl$R$QN);
    if (D == 1'b1 && GN == 1'b0 )
       (posedge  R *> (QN -: 1'b0)) = (tplh$R$QN, tphl$R$QN);
    if (D == 1'b1 && GN == 1'b1 )
       (posedge  R *> (QN -: 1'b0)) = ( tphl$R$QN);

   endspecify
endmodule //LATNRPQNX4MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATNRPQNX3MA10TR (QN, D, GN, R);
output  QN;
input  D, GN, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

not       XX0 (xRN, R);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$QN   = 1.0,
      tphl$D$QN   = 1.0,
      tplh$GN$QN   = 1.0,
      tphl$GN$QN   = 1.0,
      tplh$R$QN   = 1.0,
      tphl$R$QN   = 1.0,
      tsetup$D$GN = 1.0,
      thold$D$GN  = 0.5,
      tsetup$D$R = 1.0,
      thold$D$R  = 0.5,
      tsetup$GN$R = 1.0,
      thold$GN$R  = 0.5,
      tsetup$R$GN = 1.0,
      thold$R$GN  = 0.5,
      tminpwh$R    = 1.0,
      tminpwl$GN  = 1.0,
      tperiod$GN  = 1.0;
    // path delays
    if (SandR)
      (negedge GN *> (QN    -: D)) = (tplh$GN$QN,    tphl$GN$QN);
    if (SandRandCLK)
      ( D *> QN ) = (tplh$D$QN, tphl$D$QN );
    $setuphold(posedge GN, negedge R, tsetup$R$GN,thold$R$GN, NOTIFIER);
    $width(posedge R, tminpwh$R, 0, NOTIFIER);
    // timing checks 1
    $setuphold(posedge GN &&& (SandR == 1), posedge D, tsetup$D$GN,thold$D$GN, NOTIFIER);
    $setuphold(posedge GN &&& (SandR == 1), negedge D, tsetup$D$GN,thold$D$GN, NOTIFIER);
    $width(negedge GN &&& (SandR == 1), tminpwl$GN, 0, NOTIFIER);
    $period(posedge GN &&& (SandR == 1), tperiod$GN, NOTIFIER);
    if (D == 1'b0 && GN == 1'b1 )
       (posedge  R *> (QN -: 1'b0)) = ( tphl$R$QN);
    if (D == 1'b1 && GN == 1'b0 )
       (posedge  R *> (QN -: 1'b0)) = (tplh$R$QN, tphl$R$QN);
    if (D == 1'b1 && GN == 1'b1 )
       (posedge  R *> (QN -: 1'b0)) = ( tphl$R$QN);

   endspecify
endmodule //LATNRPQNX3MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATNRPQNX2MA10TR (QN, D, GN, R);
output  QN;
input  D, GN, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

not       XX0 (xRN, R);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$QN   = 1.0,
      tphl$D$QN   = 1.0,
      tplh$GN$QN   = 1.0,
      tphl$GN$QN   = 1.0,
      tplh$R$QN   = 1.0,
      tphl$R$QN   = 1.0,
      tsetup$D$GN = 1.0,
      thold$D$GN  = 0.5,
      tsetup$D$R = 1.0,
      thold$D$R  = 0.5,
      tsetup$GN$R = 1.0,
      thold$GN$R  = 0.5,
      tsetup$R$GN = 1.0,
      thold$R$GN  = 0.5,
      tminpwh$R    = 1.0,
      tminpwl$GN  = 1.0,
      tperiod$GN  = 1.0;
    // path delays
    if (SandR)
      (negedge GN *> (QN    -: D)) = (tplh$GN$QN,    tphl$GN$QN);
    if (SandRandCLK)
      ( D *> QN ) = (tplh$D$QN, tphl$D$QN );
    $setuphold(posedge GN, negedge R, tsetup$R$GN,thold$R$GN, NOTIFIER);
    $width(posedge R, tminpwh$R, 0, NOTIFIER);
    // timing checks 1
    $setuphold(posedge GN &&& (SandR == 1), posedge D, tsetup$D$GN,thold$D$GN, NOTIFIER);
    $setuphold(posedge GN &&& (SandR == 1), negedge D, tsetup$D$GN,thold$D$GN, NOTIFIER);
    $width(negedge GN &&& (SandR == 1), tminpwl$GN, 0, NOTIFIER);
    $period(posedge GN &&& (SandR == 1), tperiod$GN, NOTIFIER);
    if (D == 1'b0 && GN == 1'b1 )
       (posedge  R *> (QN -: 1'b0)) = ( tphl$R$QN);
    if (D == 1'b1 && GN == 1'b0 )
       (posedge  R *> (QN -: 1'b0)) = (tplh$R$QN, tphl$R$QN);
    if (D == 1'b1 && GN == 1'b1 )
       (posedge  R *> (QN -: 1'b0)) = ( tphl$R$QN);

   endspecify
endmodule //LATNRPQNX2MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATNRPQNX1MA10TR (QN, D, GN, R);
output  QN;
input  D, GN, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

not       XX0 (xRN, R);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$QN   = 1.0,
      tphl$D$QN   = 1.0,
      tplh$GN$QN   = 1.0,
      tphl$GN$QN   = 1.0,
      tplh$R$QN   = 1.0,
      tphl$R$QN   = 1.0,
      tsetup$D$GN = 1.0,
      thold$D$GN  = 0.5,
      tsetup$D$R = 1.0,
      thold$D$R  = 0.5,
      tsetup$GN$R = 1.0,
      thold$GN$R  = 0.5,
      tsetup$R$GN = 1.0,
      thold$R$GN  = 0.5,
      tminpwh$R    = 1.0,
      tminpwl$GN  = 1.0,
      tperiod$GN  = 1.0;
    // path delays
    if (SandR)
      (negedge GN *> (QN    -: D)) = (tplh$GN$QN,    tphl$GN$QN);
    if (SandRandCLK)
      ( D *> QN ) = (tplh$D$QN, tphl$D$QN );
    $setuphold(posedge GN, negedge R, tsetup$R$GN,thold$R$GN, NOTIFIER);
    $width(posedge R, tminpwh$R, 0, NOTIFIER);
    // timing checks 1
    $setuphold(posedge GN &&& (SandR == 1), posedge D, tsetup$D$GN,thold$D$GN, NOTIFIER);
    $setuphold(posedge GN &&& (SandR == 1), negedge D, tsetup$D$GN,thold$D$GN, NOTIFIER);
    $width(negedge GN &&& (SandR == 1), tminpwl$GN, 0, NOTIFIER);
    $period(posedge GN &&& (SandR == 1), tperiod$GN, NOTIFIER);
    if (D == 1'b0 && GN == 1'b1 )
       (posedge  R *> (QN -: 1'b0)) = ( tphl$R$QN);
    if (D == 1'b1 && GN == 1'b0 )
       (posedge  R *> (QN -: 1'b0)) = (tplh$R$QN, tphl$R$QN);
    if (D == 1'b1 && GN == 1'b1 )
       (posedge  R *> (QN -: 1'b0)) = ( tphl$R$QN);

   endspecify
endmodule //LATNRPQNX1MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATNRPQNX0P5MA10TR (QN, D, GN, R);
output  QN;
input  D, GN, R;
reg NOTIFIER;
supply1 xSN;
supply1 dSN;

not       XX0 (xRN, R);

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$QN   = 1.0,
      tphl$D$QN   = 1.0,
      tplh$GN$QN   = 1.0,
      tphl$GN$QN   = 1.0,
      tplh$R$QN   = 1.0,
      tphl$R$QN   = 1.0,
      tsetup$D$GN = 1.0,
      thold$D$GN  = 0.5,
      tsetup$D$R = 1.0,
      thold$D$R  = 0.5,
      tsetup$GN$R = 1.0,
      thold$GN$R  = 0.5,
      tsetup$R$GN = 1.0,
      thold$R$GN  = 0.5,
      tminpwh$R    = 1.0,
      tminpwl$GN  = 1.0,
      tperiod$GN  = 1.0;
    // path delays
    if (SandR)
      (negedge GN *> (QN    -: D)) = (tplh$GN$QN,    tphl$GN$QN);
    if (SandRandCLK)
      ( D *> QN ) = (tplh$D$QN, tphl$D$QN );
    $setuphold(posedge GN, negedge R, tsetup$R$GN,thold$R$GN, NOTIFIER);
    $width(posedge R, tminpwh$R, 0, NOTIFIER);
    // timing checks 1
    $setuphold(posedge GN &&& (SandR == 1), posedge D, tsetup$D$GN,thold$D$GN, NOTIFIER);
    $setuphold(posedge GN &&& (SandR == 1), negedge D, tsetup$D$GN,thold$D$GN, NOTIFIER);
    $width(negedge GN &&& (SandR == 1), tminpwl$GN, 0, NOTIFIER);
    $period(posedge GN &&& (SandR == 1), tperiod$GN, NOTIFIER);
    if (D == 1'b0 && GN == 1'b1 )
       (posedge  R *> (QN -: 1'b0)) = ( tphl$R$QN);
    if (D == 1'b1 && GN == 1'b0 )
       (posedge  R *> (QN -: 1'b0)) = (tplh$R$QN, tphl$R$QN);
    if (D == 1'b1 && GN == 1'b1 )
       (posedge  R *> (QN -: 1'b0)) = ( tphl$R$QN);

   endspecify
endmodule //LATNRPQNX0P5MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATNQNX4MA10TR (QN, D, GN);
output  QN;
input  D, GN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$QN   = 1.0,
      tphl$D$QN   = 1.0,
      tplh$GN$QN   = 1.0,
      tphl$GN$QN   = 1.0,
      tsetup$D$GN = 1.0,
      thold$D$GN  = 0.5,
      tminpwl$GN  = 1.0,
      tperiod$GN  = 1.0;
    // path delays
    if (SandR)
      (negedge GN *> (QN    -: D)) = (tplh$GN$QN,    tphl$GN$QN);
    if (SandRandCLK)
      ( D *> QN ) = (tplh$D$QN, tphl$D$QN );
    // timing checks 1
    $setuphold(posedge GN &&& (SandR == 1), posedge D, tsetup$D$GN,thold$D$GN, NOTIFIER);
    $setuphold(posedge GN &&& (SandR == 1), negedge D, tsetup$D$GN,thold$D$GN, NOTIFIER);
    $width(negedge GN &&& (SandR == 1), tminpwl$GN, 0, NOTIFIER);
    $period(posedge GN &&& (SandR == 1), tperiod$GN, NOTIFIER);

   endspecify
endmodule //LATNQNX4MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATNQNX3MA10TR (QN, D, GN);
output  QN;
input  D, GN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$QN   = 1.0,
      tphl$D$QN   = 1.0,
      tplh$GN$QN   = 1.0,
      tphl$GN$QN   = 1.0,
      tsetup$D$GN = 1.0,
      thold$D$GN  = 0.5,
      tminpwl$GN  = 1.0,
      tperiod$GN  = 1.0;
    // path delays
    if (SandR)
      (negedge GN *> (QN    -: D)) = (tplh$GN$QN,    tphl$GN$QN);
    if (SandRandCLK)
      ( D *> QN ) = (tplh$D$QN, tphl$D$QN );
    // timing checks 1
    $setuphold(posedge GN &&& (SandR == 1), posedge D, tsetup$D$GN,thold$D$GN, NOTIFIER);
    $setuphold(posedge GN &&& (SandR == 1), negedge D, tsetup$D$GN,thold$D$GN, NOTIFIER);
    $width(negedge GN &&& (SandR == 1), tminpwl$GN, 0, NOTIFIER);
    $period(posedge GN &&& (SandR == 1), tperiod$GN, NOTIFIER);

   endspecify
endmodule //LATNQNX3MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATNQNX2MA10TR (QN, D, GN);
output  QN;
input  D, GN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$QN   = 1.0,
      tphl$D$QN   = 1.0,
      tplh$GN$QN   = 1.0,
      tphl$GN$QN   = 1.0,
      tsetup$D$GN = 1.0,
      thold$D$GN  = 0.5,
      tminpwl$GN  = 1.0,
      tperiod$GN  = 1.0;
    // path delays
    if (SandR)
      (negedge GN *> (QN    -: D)) = (tplh$GN$QN,    tphl$GN$QN);
    if (SandRandCLK)
      ( D *> QN ) = (tplh$D$QN, tphl$D$QN );
    // timing checks 1
    $setuphold(posedge GN &&& (SandR == 1), posedge D, tsetup$D$GN,thold$D$GN, NOTIFIER);
    $setuphold(posedge GN &&& (SandR == 1), negedge D, tsetup$D$GN,thold$D$GN, NOTIFIER);
    $width(negedge GN &&& (SandR == 1), tminpwl$GN, 0, NOTIFIER);
    $period(posedge GN &&& (SandR == 1), tperiod$GN, NOTIFIER);

   endspecify
endmodule //LATNQNX2MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATNQNX1MA10TR (QN, D, GN);
output  QN;
input  D, GN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$QN   = 1.0,
      tphl$D$QN   = 1.0,
      tplh$GN$QN   = 1.0,
      tphl$GN$QN   = 1.0,
      tsetup$D$GN = 1.0,
      thold$D$GN  = 0.5,
      tminpwl$GN  = 1.0,
      tperiod$GN  = 1.0;
    // path delays
    if (SandR)
      (negedge GN *> (QN    -: D)) = (tplh$GN$QN,    tphl$GN$QN);
    if (SandRandCLK)
      ( D *> QN ) = (tplh$D$QN, tphl$D$QN );
    // timing checks 1
    $setuphold(posedge GN &&& (SandR == 1), posedge D, tsetup$D$GN,thold$D$GN, NOTIFIER);
    $setuphold(posedge GN &&& (SandR == 1), negedge D, tsetup$D$GN,thold$D$GN, NOTIFIER);
    $width(negedge GN &&& (SandR == 1), tminpwl$GN, 0, NOTIFIER);
    $period(posedge GN &&& (SandR == 1), tperiod$GN, NOTIFIER);

   endspecify
endmodule //LATNQNX1MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATNQNX0P5MA10TR (QN, D, GN);
output  QN;
input  D, GN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
not      I2 (QN, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$QN   = 1.0,
      tphl$D$QN   = 1.0,
      tplh$GN$QN   = 1.0,
      tphl$GN$QN   = 1.0,
      tsetup$D$GN = 1.0,
      thold$D$GN  = 0.5,
      tminpwl$GN  = 1.0,
      tperiod$GN  = 1.0;
    // path delays
    if (SandR)
      (negedge GN *> (QN    -: D)) = (tplh$GN$QN,    tphl$GN$QN);
    if (SandRandCLK)
      ( D *> QN ) = (tplh$D$QN, tphl$D$QN );
    // timing checks 1
    $setuphold(posedge GN &&& (SandR == 1), posedge D, tsetup$D$GN,thold$D$GN, NOTIFIER);
    $setuphold(posedge GN &&& (SandR == 1), negedge D, tsetup$D$GN,thold$D$GN, NOTIFIER);
    $width(negedge GN &&& (SandR == 1), tminpwl$GN, 0, NOTIFIER);
    $period(posedge GN &&& (SandR == 1), tperiod$GN, NOTIFIER);

   endspecify
endmodule //LATNQNX0P5MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATNQX3MA10TR (Q, D, GN);
output  Q;
input  D, GN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$Q   = 1.0,
      tphl$D$Q   = 1.0,
      tplh$GN$Q   = 1.0,
      tphl$GN$Q   = 1.0,
      tsetup$D$GN = 1.0,
      thold$D$GN  = 0.5,
      tminpwl$GN  = 1.0,
      tperiod$GN  = 1.0;
    // path delays
    if (SandR)
      (negedge GN *> (Q    +: D)) = (tplh$GN$Q,    tphl$GN$Q);
    if (SandRandCLK)
      ( D *> Q ) = (tplh$D$Q, tphl$D$Q );

    // timing checks 4
    $setuphold(posedge GN &&& (SandR == 1), posedge D, tsetup$D$GN,thold$D$GN, NOTIFIER);
    $setuphold(posedge GN &&& (SandR == 1), negedge D, tsetup$D$GN,thold$D$GN, NOTIFIER); 
    $width(negedge GN &&& (SandR == 1), tminpwl$GN, 0, NOTIFIER);
    $period(negedge GN &&& (SandR == 1), tperiod$GN, NOTIFIER);


   endspecify
endmodule //LATNQX3MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATNQX2MA10TR (Q, D, GN);
output  Q;
input  D, GN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$Q   = 1.0,
      tphl$D$Q   = 1.0,
      tplh$GN$Q   = 1.0,
      tphl$GN$Q   = 1.0,
      tsetup$D$GN = 1.0,
      thold$D$GN  = 0.5,
      tminpwl$GN  = 1.0,
      tperiod$GN  = 1.0;
    // path delays
    if (SandR)
      (negedge GN *> (Q    +: D)) = (tplh$GN$Q,    tphl$GN$Q);
    if (SandRandCLK)
      ( D *> Q ) = (tplh$D$Q, tphl$D$Q );

    // timing checks 4
    $setuphold(posedge GN &&& (SandR == 1), posedge D, tsetup$D$GN,thold$D$GN, NOTIFIER);
    $setuphold(posedge GN &&& (SandR == 1), negedge D, tsetup$D$GN,thold$D$GN, NOTIFIER); 
    $width(negedge GN &&& (SandR == 1), tminpwl$GN, 0, NOTIFIER);
    $period(negedge GN &&& (SandR == 1), tperiod$GN, NOTIFIER);


   endspecify
endmodule //LATNQX2MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATNQX1MA10TR (Q, D, GN);
output  Q;
input  D, GN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$Q   = 1.0,
      tphl$D$Q   = 1.0,
      tplh$GN$Q   = 1.0,
      tphl$GN$Q   = 1.0,
      tsetup$D$GN = 1.0,
      thold$D$GN  = 0.5,
      tminpwl$GN  = 1.0,
      tperiod$GN  = 1.0;
    // path delays
    if (SandR)
      (negedge GN *> (Q    +: D)) = (tplh$GN$Q,    tphl$GN$Q);
    if (SandRandCLK)
      ( D *> Q ) = (tplh$D$Q, tphl$D$Q );

    // timing checks 4
    $setuphold(posedge GN &&& (SandR == 1), posedge D, tsetup$D$GN,thold$D$GN, NOTIFIER);
    $setuphold(posedge GN &&& (SandR == 1), negedge D, tsetup$D$GN,thold$D$GN, NOTIFIER); 
    $width(negedge GN &&& (SandR == 1), tminpwl$GN, 0, NOTIFIER);
    $period(negedge GN &&& (SandR == 1), tperiod$GN, NOTIFIER);


   endspecify
endmodule //LATNQX1MA10TR
`endcelldefine
//$Id: tlat.genpp,v 1.9 2006/05/18 09:47:16 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module LATNQX0P5MA10TR (Q, D, GN);
output  Q;
input  D, GN;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dSN, dRN;

udp_tlat I0 (n0, D, clk, xRN, xSN, NOTIFIER);
buf      I1 (Q, n0);
buf      I3 (clk, GN);
not      I4 (flgclk, GN);
and      I5 (SandR, xSN, xRN);
and      I6 (SandRandCLK, xSN,xRN,flgclk);
 specify
   specparam 
   //timing parameters
      tplh$D$Q   = 1.0,
      tphl$D$Q   = 1.0,
      tplh$GN$Q   = 1.0,
      tphl$GN$Q   = 1.0,
      tsetup$D$GN = 1.0,
      thold$D$GN  = 0.5,
      tminpwl$GN  = 1.0,
      tperiod$GN  = 1.0;
    // path delays
    if (SandR)
      (negedge GN *> (Q    +: D)) = (tplh$GN$Q,    tphl$GN$Q);
    if (SandRandCLK)
      ( D *> Q ) = (tplh$D$Q, tphl$D$Q );

    // timing checks 4
    $setuphold(posedge GN &&& (SandR == 1), posedge D, tsetup$D$GN,thold$D$GN, NOTIFIER);
    $setuphold(posedge GN &&& (SandR == 1), negedge D, tsetup$D$GN,thold$D$GN, NOTIFIER); 
    $width(negedge GN &&& (SandR == 1), tminpwl$GN, 0, NOTIFIER);
    $period(negedge GN &&& (SandR == 1), tperiod$GN, NOTIFIER);


   endspecify
endmodule //LATNQX0P5MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX9MA10TR (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX9MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX9BA10TR (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX9BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX7P5MA10TR (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX7P5MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX7P5BA10TR (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX7P5BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX6MA10TR (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX6MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX6BA10TR (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX6BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX5MA10TR (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX5MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX5BA10TR (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX5BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX4MA10TR (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX4MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX4BA10TR (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX4BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX3P5MA10TR (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX3P5MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX3P5BA10TR (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX3P5BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX3MA10TR (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX3MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX3BA10TR (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX3BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX2P5MA10TR (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX2P5MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX2P5BA10TR (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX2P5BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX2MA10TR (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX2MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX2BA10TR (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX2BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX1P7MA10TR (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX1P7MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX1P7BA10TR (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX1P7BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX1P4MA10TR (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX1P4MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX1P4BA10TR (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX1P4BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX1P2MA10TR (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX1P2MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX1P2BA10TR (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX1P2BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX1MA10TR (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX1MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX1BA10TR (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX1BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX16MA10TR (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX16MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX16BA10TR (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX16BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX13MA10TR (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX13MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX13BA10TR (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX13BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX11MA10TR (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX11MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX11BA10TR (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX11BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX0P8MA10TR (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX0P8MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX0P8BA10TR (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX0P8BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX0P7MA10TR (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX0P7MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX0P7BA10TR (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX0P7BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX0P6MA10TR (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX0P6MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX0P6BA10TR (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX0P6BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX0P5MA10TR (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX0P5MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module INVX0P5BA10TR (Y, A);
output Y;
input A;

  not I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // INVX0P5BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module FRICGX9BA10TR (ECK, CK);
output ECK;
input CK;

  buf I0(ECK, CK);
  specify
    // delay parameters
    specparam
      tplh$CK$ECK = 1.0,
      tphl$CK$ECK = 1.0;

    // path delays
    (CK *> ECK) = (tplh$CK$ECK, tphl$CK$ECK);
  endspecify

endmodule // FRICGX9BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module FRICGX7P5BA10TR (ECK, CK);
output ECK;
input CK;

  buf I0(ECK, CK);
  specify
    // delay parameters
    specparam
      tplh$CK$ECK = 1.0,
      tphl$CK$ECK = 1.0;

    // path delays
    (CK *> ECK) = (tplh$CK$ECK, tphl$CK$ECK);
  endspecify

endmodule // FRICGX7P5BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module FRICGX6BA10TR (ECK, CK);
output ECK;
input CK;

  buf I0(ECK, CK);
  specify
    // delay parameters
    specparam
      tplh$CK$ECK = 1.0,
      tphl$CK$ECK = 1.0;

    // path delays
    (CK *> ECK) = (tplh$CK$ECK, tphl$CK$ECK);
  endspecify

endmodule // FRICGX6BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module FRICGX5BA10TR (ECK, CK);
output ECK;
input CK;

  buf I0(ECK, CK);
  specify
    // delay parameters
    specparam
      tplh$CK$ECK = 1.0,
      tphl$CK$ECK = 1.0;

    // path delays
    (CK *> ECK) = (tplh$CK$ECK, tphl$CK$ECK);
  endspecify

endmodule // FRICGX5BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module FRICGX4BA10TR (ECK, CK);
output ECK;
input CK;

  buf I0(ECK, CK);
  specify
    // delay parameters
    specparam
      tplh$CK$ECK = 1.0,
      tphl$CK$ECK = 1.0;

    // path delays
    (CK *> ECK) = (tplh$CK$ECK, tphl$CK$ECK);
  endspecify

endmodule // FRICGX4BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module FRICGX3P5BA10TR (ECK, CK);
output ECK;
input CK;

  buf I0(ECK, CK);
  specify
    // delay parameters
    specparam
      tplh$CK$ECK = 1.0,
      tphl$CK$ECK = 1.0;

    // path delays
    (CK *> ECK) = (tplh$CK$ECK, tphl$CK$ECK);
  endspecify

endmodule // FRICGX3P5BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module FRICGX3BA10TR (ECK, CK);
output ECK;
input CK;

  buf I0(ECK, CK);
  specify
    // delay parameters
    specparam
      tplh$CK$ECK = 1.0,
      tphl$CK$ECK = 1.0;

    // path delays
    (CK *> ECK) = (tplh$CK$ECK, tphl$CK$ECK);
  endspecify

endmodule // FRICGX3BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module FRICGX2P5BA10TR (ECK, CK);
output ECK;
input CK;

  buf I0(ECK, CK);
  specify
    // delay parameters
    specparam
      tplh$CK$ECK = 1.0,
      tphl$CK$ECK = 1.0;

    // path delays
    (CK *> ECK) = (tplh$CK$ECK, tphl$CK$ECK);
  endspecify

endmodule // FRICGX2P5BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module FRICGX2BA10TR (ECK, CK);
output ECK;
input CK;

  buf I0(ECK, CK);
  specify
    // delay parameters
    specparam
      tplh$CK$ECK = 1.0,
      tphl$CK$ECK = 1.0;

    // path delays
    (CK *> ECK) = (tplh$CK$ECK, tphl$CK$ECK);
  endspecify

endmodule // FRICGX2BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module FRICGX1P7BA10TR (ECK, CK);
output ECK;
input CK;

  buf I0(ECK, CK);
  specify
    // delay parameters
    specparam
      tplh$CK$ECK = 1.0,
      tphl$CK$ECK = 1.0;

    // path delays
    (CK *> ECK) = (tplh$CK$ECK, tphl$CK$ECK);
  endspecify

endmodule // FRICGX1P7BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module FRICGX1P4BA10TR (ECK, CK);
output ECK;
input CK;

  buf I0(ECK, CK);
  specify
    // delay parameters
    specparam
      tplh$CK$ECK = 1.0,
      tphl$CK$ECK = 1.0;

    // path delays
    (CK *> ECK) = (tplh$CK$ECK, tphl$CK$ECK);
  endspecify

endmodule // FRICGX1P4BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module FRICGX1P2BA10TR (ECK, CK);
output ECK;
input CK;

  buf I0(ECK, CK);
  specify
    // delay parameters
    specparam
      tplh$CK$ECK = 1.0,
      tphl$CK$ECK = 1.0;

    // path delays
    (CK *> ECK) = (tplh$CK$ECK, tphl$CK$ECK);
  endspecify

endmodule // FRICGX1P2BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module FRICGX1BA10TR (ECK, CK);
output ECK;
input CK;

  buf I0(ECK, CK);
  specify
    // delay parameters
    specparam
      tplh$CK$ECK = 1.0,
      tphl$CK$ECK = 1.0;

    // path delays
    (CK *> ECK) = (tplh$CK$ECK, tphl$CK$ECK);
  endspecify

endmodule // FRICGX1BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module FRICGX16BA10TR (ECK, CK);
output ECK;
input CK;

  buf I0(ECK, CK);
  specify
    // delay parameters
    specparam
      tplh$CK$ECK = 1.0,
      tphl$CK$ECK = 1.0;

    // path delays
    (CK *> ECK) = (tplh$CK$ECK, tphl$CK$ECK);
  endspecify

endmodule // FRICGX16BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module FRICGX13BA10TR (ECK, CK);
output ECK;
input CK;

  buf I0(ECK, CK);
  specify
    // delay parameters
    specparam
      tplh$CK$ECK = 1.0,
      tphl$CK$ECK = 1.0;

    // path delays
    (CK *> ECK) = (tplh$CK$ECK, tphl$CK$ECK);
  endspecify

endmodule // FRICGX13BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module FRICGX11BA10TR (ECK, CK);
output ECK;
input CK;

  buf I0(ECK, CK);
  specify
    // delay parameters
    specparam
      tplh$CK$ECK = 1.0,
      tphl$CK$ECK = 1.0;

    // path delays
    (CK *> ECK) = (tplh$CK$ECK, tphl$CK$ECK);
  endspecify

endmodule // FRICGX11BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module FRICGX0P8BA10TR (ECK, CK);
output ECK;
input CK;

  buf I0(ECK, CK);
  specify
    // delay parameters
    specparam
      tplh$CK$ECK = 1.0,
      tphl$CK$ECK = 1.0;

    // path delays
    (CK *> ECK) = (tplh$CK$ECK, tphl$CK$ECK);
  endspecify

endmodule // FRICGX0P8BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module FRICGX0P7BA10TR (ECK, CK);
output ECK;
input CK;

  buf I0(ECK, CK);
  specify
    // delay parameters
    specparam
      tplh$CK$ECK = 1.0,
      tphl$CK$ECK = 1.0;

    // path delays
    (CK *> ECK) = (tplh$CK$ECK, tphl$CK$ECK);
  endspecify

endmodule // FRICGX0P7BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module FRICGX0P6BA10TR (ECK, CK);
output ECK;
input CK;

  buf I0(ECK, CK);
  specify
    // delay parameters
    specparam
      tplh$CK$ECK = 1.0,
      tphl$CK$ECK = 1.0;

    // path delays
    (CK *> ECK) = (tplh$CK$ECK, tphl$CK$ECK);
  endspecify

endmodule // FRICGX0P6BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module FRICGX0P5BA10TR (ECK, CK);
output ECK;
input CK;

  buf I0(ECK, CK);
  specify
    // delay parameters
    specparam
      tplh$CK$ECK = 1.0,
      tphl$CK$ECK = 1.0;

    // path delays
    (CK *> ECK) = (tplh$CK$ECK, tphl$CK$ECK);
  endspecify

endmodule // FRICGX0P5BA10TR
`endcelldefine
//$Id: edff.genpp,v 1.12 2006/07/19 10:36:43 rmouli Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module ESDFFQNX3MA10TR (QN, D, CK, E, SE, SI);
output QN;
input D, CK, E, SE, SI;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff I0 (n0, D, CK, xRN, SI, SE, E, NOTIFIER);
   not       I1 (QN, n0);
   and       I3 (SandR, xSN, xRN);
   buf       I4 (scan, SE);
   not       I5 (notscan, SE);
   and       I6 (Dcheck, notscan, E);
  specify
    specparam 
      tplh$CK$QN    = 1.0,
      tphl$CK$QN    = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK  = 0.5,
      tsetup$CK$CK = 1.0,
      thold$CK$CK  = 0.5,
      tsetup$E$CK = 1.0,
      thold$E$CK  = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK  = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK  = 0.5,
      
      tminpwl$CK  = 1.0,
      tminpwh$CK  = 1.0,
      tperiod$CK  = 1.0;
    // path delays
     if (scan)
	(posedge CK *> (QN    -: SI)) = (tplh$CK$QN,    tphl$CK$QN);
     if (notscan)
	(posedge CK *> (QN    -: E)) = (tplh$CK$QN,    tphl$CK$QN);
     if (Dcheck)
	(posedge CK *> (QN    -: D)) = (tplh$CK$QN,    tphl$CK$QN);
     (posedge CK *> (QN    -: SE)) = (tplh$CK$QN,    tphl$CK$QN);
     // timing checks
     $setuphold(posedge CK &&& (Dcheck == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
     $setuphold(posedge CK &&& (Dcheck == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
     $setuphold(posedge CK &&& (scan == 1), posedge SI, tsetup$SI$CK ,thold$SI$CK, NOTIFIER);
     $setuphold(posedge CK &&& (scan == 1), negedge SI, tsetup$SI$CK ,thold$SI$CK, NOTIFIER);
     $setuphold(posedge CK &&& (notscan == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
     $setuphold(posedge CK &&& (notscan == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
     $setuphold(posedge CK, posedge SE,  tsetup$SE$CK ,thold$SE$CK , NOTIFIER);
     $setuphold(posedge CK, negedge SE,  tsetup$SE$CK ,thold$SE$CK , NOTIFIER);
     $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
     $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
     $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
  endspecify
endmodule // ESDFFQNX3MA10TR
`endcelldefine


//$Id: edff.genpp,v 1.12 2006/07/19 10:36:43 rmouli Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module ESDFFQNX2MA10TR (QN, D, CK, E, SE, SI);
output QN;
input D, CK, E, SE, SI;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff I0 (n0, D, CK, xRN, SI, SE, E, NOTIFIER);
   not       I1 (QN, n0);
   and       I3 (SandR, xSN, xRN);
   buf       I4 (scan, SE);
   not       I5 (notscan, SE);
   and       I6 (Dcheck, notscan, E);
  specify
    specparam 
      tplh$CK$QN    = 1.0,
      tphl$CK$QN    = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK  = 0.5,
      tsetup$CK$CK = 1.0,
      thold$CK$CK  = 0.5,
      tsetup$E$CK = 1.0,
      thold$E$CK  = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK  = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK  = 0.5,
      
      tminpwl$CK  = 1.0,
      tminpwh$CK  = 1.0,
      tperiod$CK  = 1.0;
    // path delays
     if (scan)
	(posedge CK *> (QN    -: SI)) = (tplh$CK$QN,    tphl$CK$QN);
     if (notscan)
	(posedge CK *> (QN    -: E)) = (tplh$CK$QN,    tphl$CK$QN);
     if (Dcheck)
	(posedge CK *> (QN    -: D)) = (tplh$CK$QN,    tphl$CK$QN);
     (posedge CK *> (QN    -: SE)) = (tplh$CK$QN,    tphl$CK$QN);
     // timing checks
     $setuphold(posedge CK &&& (Dcheck == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
     $setuphold(posedge CK &&& (Dcheck == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
     $setuphold(posedge CK &&& (scan == 1), posedge SI, tsetup$SI$CK ,thold$SI$CK, NOTIFIER);
     $setuphold(posedge CK &&& (scan == 1), negedge SI, tsetup$SI$CK ,thold$SI$CK, NOTIFIER);
     $setuphold(posedge CK &&& (notscan == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
     $setuphold(posedge CK &&& (notscan == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
     $setuphold(posedge CK, posedge SE,  tsetup$SE$CK ,thold$SE$CK , NOTIFIER);
     $setuphold(posedge CK, negedge SE,  tsetup$SE$CK ,thold$SE$CK , NOTIFIER);
     $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
     $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
     $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
  endspecify
endmodule // ESDFFQNX2MA10TR
`endcelldefine


//$Id: edff.genpp,v 1.12 2006/07/19 10:36:43 rmouli Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module ESDFFQNX1MA10TR (QN, D, CK, E, SE, SI);
output QN;
input D, CK, E, SE, SI;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff I0 (n0, D, CK, xRN, SI, SE, E, NOTIFIER);
   not       I1 (QN, n0);
   and       I3 (SandR, xSN, xRN);
   buf       I4 (scan, SE);
   not       I5 (notscan, SE);
   and       I6 (Dcheck, notscan, E);
  specify
    specparam 
      tplh$CK$QN    = 1.0,
      tphl$CK$QN    = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK  = 0.5,
      tsetup$CK$CK = 1.0,
      thold$CK$CK  = 0.5,
      tsetup$E$CK = 1.0,
      thold$E$CK  = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK  = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK  = 0.5,
      
      tminpwl$CK  = 1.0,
      tminpwh$CK  = 1.0,
      tperiod$CK  = 1.0;
    // path delays
     if (scan)
	(posedge CK *> (QN    -: SI)) = (tplh$CK$QN,    tphl$CK$QN);
     if (notscan)
	(posedge CK *> (QN    -: E)) = (tplh$CK$QN,    tphl$CK$QN);
     if (Dcheck)
	(posedge CK *> (QN    -: D)) = (tplh$CK$QN,    tphl$CK$QN);
     (posedge CK *> (QN    -: SE)) = (tplh$CK$QN,    tphl$CK$QN);
     // timing checks
     $setuphold(posedge CK &&& (Dcheck == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
     $setuphold(posedge CK &&& (Dcheck == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
     $setuphold(posedge CK &&& (scan == 1), posedge SI, tsetup$SI$CK ,thold$SI$CK, NOTIFIER);
     $setuphold(posedge CK &&& (scan == 1), negedge SI, tsetup$SI$CK ,thold$SI$CK, NOTIFIER);
     $setuphold(posedge CK &&& (notscan == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
     $setuphold(posedge CK &&& (notscan == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
     $setuphold(posedge CK, posedge SE,  tsetup$SE$CK ,thold$SE$CK , NOTIFIER);
     $setuphold(posedge CK, negedge SE,  tsetup$SE$CK ,thold$SE$CK , NOTIFIER);
     $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
     $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
     $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
  endspecify
endmodule // ESDFFQNX1MA10TR
`endcelldefine


//$Id: edff.genpp,v 1.12 2006/07/19 10:36:43 rmouli Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module ESDFFQNX0P5MA10TR (QN, D, CK, E, SE, SI);
output QN;
input D, CK, E, SE, SI;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff I0 (n0, D, CK, xRN, SI, SE, E, NOTIFIER);
   not       I1 (QN, n0);
   and       I3 (SandR, xSN, xRN);
   buf       I4 (scan, SE);
   not       I5 (notscan, SE);
   and       I6 (Dcheck, notscan, E);
  specify
    specparam 
      tplh$CK$QN    = 1.0,
      tphl$CK$QN    = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK  = 0.5,
      tsetup$CK$CK = 1.0,
      thold$CK$CK  = 0.5,
      tsetup$E$CK = 1.0,
      thold$E$CK  = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK  = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK  = 0.5,
      
      tminpwl$CK  = 1.0,
      tminpwh$CK  = 1.0,
      tperiod$CK  = 1.0;
    // path delays
     if (scan)
	(posedge CK *> (QN    -: SI)) = (tplh$CK$QN,    tphl$CK$QN);
     if (notscan)
	(posedge CK *> (QN    -: E)) = (tplh$CK$QN,    tphl$CK$QN);
     if (Dcheck)
	(posedge CK *> (QN    -: D)) = (tplh$CK$QN,    tphl$CK$QN);
     (posedge CK *> (QN    -: SE)) = (tplh$CK$QN,    tphl$CK$QN);
     // timing checks
     $setuphold(posedge CK &&& (Dcheck == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
     $setuphold(posedge CK &&& (Dcheck == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
     $setuphold(posedge CK &&& (scan == 1), posedge SI, tsetup$SI$CK ,thold$SI$CK, NOTIFIER);
     $setuphold(posedge CK &&& (scan == 1), negedge SI, tsetup$SI$CK ,thold$SI$CK, NOTIFIER);
     $setuphold(posedge CK &&& (notscan == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
     $setuphold(posedge CK &&& (notscan == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
     $setuphold(posedge CK, posedge SE,  tsetup$SE$CK ,thold$SE$CK , NOTIFIER);
     $setuphold(posedge CK, negedge SE,  tsetup$SE$CK ,thold$SE$CK , NOTIFIER);
     $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
     $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
     $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
  endspecify
endmodule // ESDFFQNX0P5MA10TR
`endcelldefine


//$Id: edff.genpp,v 1.12 2006/07/19 10:36:43 rmouli Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module ESDFFQX3MA10TR (Q, D, CK, E, SE, SI);
output Q;
input D, CK, E, SE, SI;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff I0 (n0, D, CK, xRN, SI, SE, E, NOTIFIER);
   buf       I1 (Q, n0);
   and       I3 (SandR, xSN, xRN);
   buf       I4 (scan, SE);
   not       I5 (notscan, SE);
   and       I6 (Dcheck, notscan, E);
  specify
    specparam 
      tplh$CK$Q    = 1.0,
      tphl$CK$Q    = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK  = 0.5,
      tsetup$CK$CK = 1.0,
      thold$CK$CK  = 0.5,
      tsetup$E$CK = 1.0,
      thold$E$CK  = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK  = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK  = 0.5,
      
      tminpwl$CK  = 1.0,
      tminpwh$CK  = 1.0,
      tperiod$CK  = 1.0;
    // path delays
     if (scan)
	(posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);
     if (notscan)
	(posedge CK *> (Q    +: E)) = (tplh$CK$Q,    tphl$CK$Q);
     if (Dcheck)
	(posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
     (posedge CK *> (Q    +: SE)) = (tplh$CK$Q,    tphl$CK$Q);
     // timing checks
     $setuphold(posedge CK &&& (Dcheck == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
     $setuphold(posedge CK &&& (Dcheck == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
     $setuphold(posedge CK &&& (scan == 1), posedge SI, tsetup$SI$CK ,thold$SI$CK, NOTIFIER);
     $setuphold(posedge CK &&& (scan == 1), negedge SI, tsetup$SI$CK ,thold$SI$CK, NOTIFIER);
     $setuphold(posedge CK &&& (notscan == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
     $setuphold(posedge CK &&& (notscan == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
     $setuphold(posedge CK, posedge SE,  tsetup$SE$CK ,thold$SE$CK , NOTIFIER);
     $setuphold(posedge CK, negedge SE,  tsetup$SE$CK ,thold$SE$CK , NOTIFIER);
     $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
     $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
     $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
  endspecify
endmodule // ESDFFQX3MA10TR
`endcelldefine


//$Id: edff.genpp,v 1.12 2006/07/19 10:36:43 rmouli Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module ESDFFQX2MA10TR (Q, D, CK, E, SE, SI);
output Q;
input D, CK, E, SE, SI;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff I0 (n0, D, CK, xRN, SI, SE, E, NOTIFIER);
   buf       I1 (Q, n0);
   and       I3 (SandR, xSN, xRN);
   buf       I4 (scan, SE);
   not       I5 (notscan, SE);
   and       I6 (Dcheck, notscan, E);
  specify
    specparam 
      tplh$CK$Q    = 1.0,
      tphl$CK$Q    = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK  = 0.5,
      tsetup$CK$CK = 1.0,
      thold$CK$CK  = 0.5,
      tsetup$E$CK = 1.0,
      thold$E$CK  = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK  = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK  = 0.5,
      
      tminpwl$CK  = 1.0,
      tminpwh$CK  = 1.0,
      tperiod$CK  = 1.0;
    // path delays
     if (scan)
	(posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);
     if (notscan)
	(posedge CK *> (Q    +: E)) = (tplh$CK$Q,    tphl$CK$Q);
     if (Dcheck)
	(posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
     (posedge CK *> (Q    +: SE)) = (tplh$CK$Q,    tphl$CK$Q);
     // timing checks
     $setuphold(posedge CK &&& (Dcheck == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
     $setuphold(posedge CK &&& (Dcheck == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
     $setuphold(posedge CK &&& (scan == 1), posedge SI, tsetup$SI$CK ,thold$SI$CK, NOTIFIER);
     $setuphold(posedge CK &&& (scan == 1), negedge SI, tsetup$SI$CK ,thold$SI$CK, NOTIFIER);
     $setuphold(posedge CK &&& (notscan == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
     $setuphold(posedge CK &&& (notscan == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
     $setuphold(posedge CK, posedge SE,  tsetup$SE$CK ,thold$SE$CK , NOTIFIER);
     $setuphold(posedge CK, negedge SE,  tsetup$SE$CK ,thold$SE$CK , NOTIFIER);
     $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
     $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
     $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
  endspecify
endmodule // ESDFFQX2MA10TR
`endcelldefine


//$Id: edff.genpp,v 1.12 2006/07/19 10:36:43 rmouli Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module ESDFFQX1MA10TR (Q, D, CK, E, SE, SI);
output Q;
input D, CK, E, SE, SI;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff I0 (n0, D, CK, xRN, SI, SE, E, NOTIFIER);
   buf       I1 (Q, n0);
   and       I3 (SandR, xSN, xRN);
   buf       I4 (scan, SE);
   not       I5 (notscan, SE);
   and       I6 (Dcheck, notscan, E);
  specify
    specparam 
      tplh$CK$Q    = 1.0,
      tphl$CK$Q    = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK  = 0.5,
      tsetup$CK$CK = 1.0,
      thold$CK$CK  = 0.5,
      tsetup$E$CK = 1.0,
      thold$E$CK  = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK  = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK  = 0.5,
      
      tminpwl$CK  = 1.0,
      tminpwh$CK  = 1.0,
      tperiod$CK  = 1.0;
    // path delays
     if (scan)
	(posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);
     if (notscan)
	(posedge CK *> (Q    +: E)) = (tplh$CK$Q,    tphl$CK$Q);
     if (Dcheck)
	(posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
     (posedge CK *> (Q    +: SE)) = (tplh$CK$Q,    tphl$CK$Q);
     // timing checks
     $setuphold(posedge CK &&& (Dcheck == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
     $setuphold(posedge CK &&& (Dcheck == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
     $setuphold(posedge CK &&& (scan == 1), posedge SI, tsetup$SI$CK ,thold$SI$CK, NOTIFIER);
     $setuphold(posedge CK &&& (scan == 1), negedge SI, tsetup$SI$CK ,thold$SI$CK, NOTIFIER);
     $setuphold(posedge CK &&& (notscan == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
     $setuphold(posedge CK &&& (notscan == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
     $setuphold(posedge CK, posedge SE,  tsetup$SE$CK ,thold$SE$CK , NOTIFIER);
     $setuphold(posedge CK, negedge SE,  tsetup$SE$CK ,thold$SE$CK , NOTIFIER);
     $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
     $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
     $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
  endspecify
endmodule // ESDFFQX1MA10TR
`endcelldefine


//$Id: edff.genpp,v 1.12 2006/07/19 10:36:43 rmouli Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module ESDFFQX0P5MA10TR (Q, D, CK, E, SE, SI);
output Q;
input D, CK, E, SE, SI;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

   udp_sedff I0 (n0, D, CK, xRN, SI, SE, E, NOTIFIER);
   buf       I1 (Q, n0);
   and       I3 (SandR, xSN, xRN);
   buf       I4 (scan, SE);
   not       I5 (notscan, SE);
   and       I6 (Dcheck, notscan, E);
  specify
    specparam 
      tplh$CK$Q    = 1.0,
      tphl$CK$Q    = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK  = 0.5,
      tsetup$CK$CK = 1.0,
      thold$CK$CK  = 0.5,
      tsetup$E$CK = 1.0,
      thold$E$CK  = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK  = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK  = 0.5,
      
      tminpwl$CK  = 1.0,
      tminpwh$CK  = 1.0,
      tperiod$CK  = 1.0;
    // path delays
     if (scan)
	(posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);
     if (notscan)
	(posedge CK *> (Q    +: E)) = (tplh$CK$Q,    tphl$CK$Q);
     if (Dcheck)
	(posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
     (posedge CK *> (Q    +: SE)) = (tplh$CK$Q,    tphl$CK$Q);
     // timing checks
     $setuphold(posedge CK &&& (Dcheck == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
     $setuphold(posedge CK &&& (Dcheck == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
     $setuphold(posedge CK &&& (scan == 1), posedge SI, tsetup$SI$CK ,thold$SI$CK, NOTIFIER);
     $setuphold(posedge CK &&& (scan == 1), negedge SI, tsetup$SI$CK ,thold$SI$CK, NOTIFIER);
     $setuphold(posedge CK &&& (notscan == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
     $setuphold(posedge CK &&& (notscan == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
     $setuphold(posedge CK, posedge SE,  tsetup$SE$CK ,thold$SE$CK , NOTIFIER);
     $setuphold(posedge CK, negedge SE,  tsetup$SE$CK ,thold$SE$CK , NOTIFIER);
     $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
     $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
     $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);
  endspecify
endmodule // ESDFFQX0P5MA10TR
`endcelldefine


//$Id: edff.genpp,v 1.12 2006/07/19 10:36:43 rmouli Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module EDFFQNX3MA10TR (QN, D, CK, E);
output QN;
input D, CK, E;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

  udp_edff I0 (n0, D, CK, xRN, xSN, E, NOTIFIER);
  not      I1 (QN, n0);
  and      I2 (flag, xRN, xSN);
  and      I3 (Dcheck, xSN, xRN, E);
  specify
    specparam 
      tplh$CK$QN    = 1.0,
      tphl$CK$QN    = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK  = 0.5,
      tsetup$CK$CK = 1.0,
      thold$CK$CK  = 0.5,
      tsetup$E$CK = 1.0,
      thold$E$CK  = 0.5,
      tminpwl$CK  = 1.0,
      tminpwh$CK  = 1.0,
      tperiod$CK  = 1.0;
    // path delays
     if (Dcheck)
        (posedge CK *> (QN -: D)) = (tplh$CK$QN, tphl$CK$QN);
     // timing checks
    $setuphold(posedge CK &&& (Dcheck == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (Dcheck == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
     $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
     $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER);
     $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
  endspecify
endmodule // EDFFQNX3MA10TR
`endcelldefine


//$Id: edff.genpp,v 1.12 2006/07/19 10:36:43 rmouli Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module EDFFQNX2MA10TR (QN, D, CK, E);
output QN;
input D, CK, E;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

  udp_edff I0 (n0, D, CK, xRN, xSN, E, NOTIFIER);
  not      I1 (QN, n0);
  and      I2 (flag, xRN, xSN);
  and      I3 (Dcheck, xSN, xRN, E);
  specify
    specparam 
      tplh$CK$QN    = 1.0,
      tphl$CK$QN    = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK  = 0.5,
      tsetup$CK$CK = 1.0,
      thold$CK$CK  = 0.5,
      tsetup$E$CK = 1.0,
      thold$E$CK  = 0.5,
      tminpwl$CK  = 1.0,
      tminpwh$CK  = 1.0,
      tperiod$CK  = 1.0;
    // path delays
     if (Dcheck)
        (posedge CK *> (QN -: D)) = (tplh$CK$QN, tphl$CK$QN);
     // timing checks
    $setuphold(posedge CK &&& (Dcheck == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (Dcheck == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
     $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
     $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER);
     $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
  endspecify
endmodule // EDFFQNX2MA10TR
`endcelldefine


//$Id: edff.genpp,v 1.12 2006/07/19 10:36:43 rmouli Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module EDFFQNX1MA10TR (QN, D, CK, E);
output QN;
input D, CK, E;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

  udp_edff I0 (n0, D, CK, xRN, xSN, E, NOTIFIER);
  not      I1 (QN, n0);
  and      I2 (flag, xRN, xSN);
  and      I3 (Dcheck, xSN, xRN, E);
  specify
    specparam 
      tplh$CK$QN    = 1.0,
      tphl$CK$QN    = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK  = 0.5,
      tsetup$CK$CK = 1.0,
      thold$CK$CK  = 0.5,
      tsetup$E$CK = 1.0,
      thold$E$CK  = 0.5,
      tminpwl$CK  = 1.0,
      tminpwh$CK  = 1.0,
      tperiod$CK  = 1.0;
    // path delays
     if (Dcheck)
        (posedge CK *> (QN -: D)) = (tplh$CK$QN, tphl$CK$QN);
     // timing checks
    $setuphold(posedge CK &&& (Dcheck == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (Dcheck == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
     $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
     $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER);
     $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
  endspecify
endmodule // EDFFQNX1MA10TR
`endcelldefine


//$Id: edff.genpp,v 1.12 2006/07/19 10:36:43 rmouli Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module EDFFQNX0P5MA10TR (QN, D, CK, E);
output QN;
input D, CK, E;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

  udp_edff I0 (n0, D, CK, xRN, xSN, E, NOTIFIER);
  not      I1 (QN, n0);
  and      I2 (flag, xRN, xSN);
  and      I3 (Dcheck, xSN, xRN, E);
  specify
    specparam 
      tplh$CK$QN    = 1.0,
      tphl$CK$QN    = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK  = 0.5,
      tsetup$CK$CK = 1.0,
      thold$CK$CK  = 0.5,
      tsetup$E$CK = 1.0,
      thold$E$CK  = 0.5,
      tminpwl$CK  = 1.0,
      tminpwh$CK  = 1.0,
      tperiod$CK  = 1.0;
    // path delays
     if (Dcheck)
        (posedge CK *> (QN -: D)) = (tplh$CK$QN, tphl$CK$QN);
     // timing checks
    $setuphold(posedge CK &&& (Dcheck == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (Dcheck == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
     $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
     $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER);
     $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
  endspecify
endmodule // EDFFQNX0P5MA10TR
`endcelldefine


//$Id: edff.genpp,v 1.12 2006/07/19 10:36:43 rmouli Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module EDFFQX3MA10TR (Q, D, CK, E);
output Q;
input D, CK, E;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

  udp_edff I0 (n0, D, CK, xRN, xSN, E, NOTIFIER);
  buf     B1 (Q, n0);
  and      I2 (flag, xRN, xSN);
  and      I3 (Dcheck, xSN, xRN, E);
  specify
    specparam 
      tplh$CK$Q    = 1.0,
      tphl$CK$Q    = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK  = 0.5,
      tsetup$CK$CK = 1.0,
      thold$CK$CK  = 0.5,
      tsetup$E$CK = 1.0,
      thold$E$CK  = 0.5,
      tminpwl$CK  = 1.0,
      tminpwh$CK  = 1.0,
      tperiod$CK  = 1.0;
    // path delays
     if (Dcheck)
        (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
     // timing checks
    $setuphold(posedge CK &&& (Dcheck == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (Dcheck == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
     $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
     $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER);
     $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
  endspecify
endmodule // EDFFQX3MA10TR
`endcelldefine


//$Id: edff.genpp,v 1.12 2006/07/19 10:36:43 rmouli Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module EDFFQX2MA10TR (Q, D, CK, E);
output Q;
input D, CK, E;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

  udp_edff I0 (n0, D, CK, xRN, xSN, E, NOTIFIER);
  buf     B1 (Q, n0);
  and      I2 (flag, xRN, xSN);
  and      I3 (Dcheck, xSN, xRN, E);
  specify
    specparam 
      tplh$CK$Q    = 1.0,
      tphl$CK$Q    = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK  = 0.5,
      tsetup$CK$CK = 1.0,
      thold$CK$CK  = 0.5,
      tsetup$E$CK = 1.0,
      thold$E$CK  = 0.5,
      tminpwl$CK  = 1.0,
      tminpwh$CK  = 1.0,
      tperiod$CK  = 1.0;
    // path delays
     if (Dcheck)
        (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
     // timing checks
    $setuphold(posedge CK &&& (Dcheck == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (Dcheck == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
     $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
     $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER);
     $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
  endspecify
endmodule // EDFFQX2MA10TR
`endcelldefine


//$Id: edff.genpp,v 1.12 2006/07/19 10:36:43 rmouli Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module EDFFQX1MA10TR (Q, D, CK, E);
output Q;
input D, CK, E;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

  udp_edff I0 (n0, D, CK, xRN, xSN, E, NOTIFIER);
  buf     B1 (Q, n0);
  and      I2 (flag, xRN, xSN);
  and      I3 (Dcheck, xSN, xRN, E);
  specify
    specparam 
      tplh$CK$Q    = 1.0,
      tphl$CK$Q    = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK  = 0.5,
      tsetup$CK$CK = 1.0,
      thold$CK$CK  = 0.5,
      tsetup$E$CK = 1.0,
      thold$E$CK  = 0.5,
      tminpwl$CK  = 1.0,
      tminpwh$CK  = 1.0,
      tperiod$CK  = 1.0;
    // path delays
     if (Dcheck)
        (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
     // timing checks
    $setuphold(posedge CK &&& (Dcheck == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (Dcheck == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
     $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
     $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER);
     $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
  endspecify
endmodule // EDFFQX1MA10TR
`endcelldefine


//$Id: edff.genpp,v 1.12 2006/07/19 10:36:43 rmouli Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module EDFFQX0P5MA10TR (Q, D, CK, E);
output Q;
input D, CK, E;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;

  udp_edff I0 (n0, D, CK, xRN, xSN, E, NOTIFIER);
  buf     B1 (Q, n0);
  and      I2 (flag, xRN, xSN);
  and      I3 (Dcheck, xSN, xRN, E);
  specify
    specparam 
      tplh$CK$Q    = 1.0,
      tphl$CK$Q    = 1.0,
      tsetup$D$CK = 1.0,
      thold$D$CK  = 0.5,
      tsetup$CK$CK = 1.0,
      thold$CK$CK  = 0.5,
      tsetup$E$CK = 1.0,
      thold$E$CK  = 0.5,
      tminpwl$CK  = 1.0,
      tminpwh$CK  = 1.0,
      tperiod$CK  = 1.0;
    // path delays
     if (Dcheck)
        (posedge CK *> (Q    +: D)) = (tplh$CK$Q,    tphl$CK$Q);
     // timing checks
    $setuphold(posedge CK &&& (Dcheck == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (Dcheck == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), posedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge E, tsetup$E$CK, thold$E$CK, NOTIFIER);
     $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
     $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER);
     $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
  endspecify
endmodule // EDFFQX0P5MA10TR
`endcelldefine


//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DLY4X0P5MA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // DLY4X0P5MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DLY2X0P5MA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // DLY2X0P5MA10TR
`endcelldefine
//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFYQX4MA10TR (Q, D, CK);
output Q;
input  D, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // DFFYQX4MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFYQX3MA10TR (Q, D, CK);
output Q;
input  D, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // DFFYQX3MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFYQX2MA10TR (Q, D, CK);
output Q;
input  D, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // DFFYQX2MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFYQX1MA10TR (Q, D, CK);
output Q;
input  D, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // DFFYQX1MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFSRPQX4MA10TR (Q, D, CK, SN, R);
output Q;
input  D, CK, SN, R;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  not   XX1 (xRN, R);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$SN$Q  = 1.0,
    tphl$SN$Q  = 1.0,
    tplh$R$Q  = 1.0,
    tphl$R$Q  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tsetup$SN$CK    = 1.0,
    thold$SN$CK    = 0.5,
    tminpwl$SN     = 1.0,
    tminpwh$SN     = 1.0,
    tsetup$R$CK    = 1.0,
    thold$R$CK    = 0.5,
    tminpwl$R     = 1.0,
    tminpwh$R     = 1.0,
    thold$R$SN = 1.0,
    thold$SN$R = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK, negedge R &&& (SN == 1'b1), tsetup$R$CK, thold$R$CK, NOTIFIER);
    $width(posedge R &&& (SN == 1'b1), tminpwh$R, 0, NOTIFIER);
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK, thold$SN$CK, NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    $hold(negedge R, negedge SN, thold$SN$R, NOTIFIER);    
    $hold(posedge SN, posedge R, thold$R$SN, NOTIFIER);    
    if (D == 1'b0 && SN == 1'b1 && CK == 1'b0)
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b0 && R == 1'b0 && CK == 1'b0)
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q); 
    if (D == 1'b0 && SN == 1'b1 && CK == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b0 && R == 1'b0 && CK == 1'b1)
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q); 
    if (D == 1'b1 && SN == 1'b1 && CK == 1'b0)
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b1 && R == 1'b0 && CK == 1'b0)
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q); 
    if (D == 1'b1 && SN == 1'b1 && CK == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b1 && R == 1'b0 && CK == 1'b1)
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q); 

   endspecify
endmodule // DFFSRPQX4MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFSRPQX3MA10TR (Q, D, CK, SN, R);
output Q;
input  D, CK, SN, R;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  not   XX1 (xRN, R);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$SN$Q  = 1.0,
    tphl$SN$Q  = 1.0,
    tplh$R$Q  = 1.0,
    tphl$R$Q  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tsetup$SN$CK    = 1.0,
    thold$SN$CK    = 0.5,
    tminpwl$SN     = 1.0,
    tminpwh$SN     = 1.0,
    tsetup$R$CK    = 1.0,
    thold$R$CK    = 0.5,
    tminpwl$R     = 1.0,
    tminpwh$R     = 1.0,
    thold$R$SN = 1.0,
    thold$SN$R = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK, negedge R &&& (SN == 1'b1), tsetup$R$CK, thold$R$CK, NOTIFIER);
    $width(posedge R &&& (SN == 1'b1), tminpwh$R, 0, NOTIFIER);
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK, thold$SN$CK, NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    $hold(negedge R, negedge SN, thold$SN$R, NOTIFIER);    
    $hold(posedge SN, posedge R, thold$R$SN, NOTIFIER);    
    if (D == 1'b0 && SN == 1'b1 && CK == 1'b0)
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b0 && R == 1'b0 && CK == 1'b0)
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q); 
    if (D == 1'b0 && SN == 1'b1 && CK == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b0 && R == 1'b0 && CK == 1'b1)
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q); 
    if (D == 1'b1 && SN == 1'b1 && CK == 1'b0)
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b1 && R == 1'b0 && CK == 1'b0)
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q); 
    if (D == 1'b1 && SN == 1'b1 && CK == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b1 && R == 1'b0 && CK == 1'b1)
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q); 

   endspecify
endmodule // DFFSRPQX3MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFSRPQX2MA10TR (Q, D, CK, SN, R);
output Q;
input  D, CK, SN, R;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  not   XX1 (xRN, R);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$SN$Q  = 1.0,
    tphl$SN$Q  = 1.0,
    tplh$R$Q  = 1.0,
    tphl$R$Q  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tsetup$SN$CK    = 1.0,
    thold$SN$CK    = 0.5,
    tminpwl$SN     = 1.0,
    tminpwh$SN     = 1.0,
    tsetup$R$CK    = 1.0,
    thold$R$CK    = 0.5,
    tminpwl$R     = 1.0,
    tminpwh$R     = 1.0,
    thold$R$SN = 1.0,
    thold$SN$R = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK, negedge R &&& (SN == 1'b1), tsetup$R$CK, thold$R$CK, NOTIFIER);
    $width(posedge R &&& (SN == 1'b1), tminpwh$R, 0, NOTIFIER);
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK, thold$SN$CK, NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    $hold(negedge R, negedge SN, thold$SN$R, NOTIFIER);    
    $hold(posedge SN, posedge R, thold$R$SN, NOTIFIER);    
    if (D == 1'b0 && SN == 1'b1 && CK == 1'b0)
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b0 && R == 1'b0 && CK == 1'b0)
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q); 
    if (D == 1'b0 && SN == 1'b1 && CK == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b0 && R == 1'b0 && CK == 1'b1)
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q); 
    if (D == 1'b1 && SN == 1'b1 && CK == 1'b0)
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b1 && R == 1'b0 && CK == 1'b0)
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q); 
    if (D == 1'b1 && SN == 1'b1 && CK == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b1 && R == 1'b0 && CK == 1'b1)
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q); 

   endspecify
endmodule // DFFSRPQX2MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFSRPQX1MA10TR (Q, D, CK, SN, R);
output Q;
input  D, CK, SN, R;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  not   XX1 (xRN, R);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$SN$Q  = 1.0,
    tphl$SN$Q  = 1.0,
    tplh$R$Q  = 1.0,
    tphl$R$Q  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tsetup$SN$CK    = 1.0,
    thold$SN$CK    = 0.5,
    tminpwl$SN     = 1.0,
    tminpwh$SN     = 1.0,
    tsetup$R$CK    = 1.0,
    thold$R$CK    = 0.5,
    tminpwl$R     = 1.0,
    tminpwh$R     = 1.0,
    thold$R$SN = 1.0,
    thold$SN$R = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK, negedge R &&& (SN == 1'b1), tsetup$R$CK, thold$R$CK, NOTIFIER);
    $width(posedge R &&& (SN == 1'b1), tminpwh$R, 0, NOTIFIER);
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK, thold$SN$CK, NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    $hold(negedge R, negedge SN, thold$SN$R, NOTIFIER);    
    $hold(posedge SN, posedge R, thold$R$SN, NOTIFIER);    
    if (D == 1'b0 && SN == 1'b1 && CK == 1'b0)
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b0 && R == 1'b0 && CK == 1'b0)
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q); 
    if (D == 1'b0 && SN == 1'b1 && CK == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b0 && R == 1'b0 && CK == 1'b1)
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q); 
    if (D == 1'b1 && SN == 1'b1 && CK == 1'b0)
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b1 && R == 1'b0 && CK == 1'b0)
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q); 
    if (D == 1'b1 && SN == 1'b1 && CK == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b1 && R == 1'b0 && CK == 1'b1)
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q); 

   endspecify
endmodule // DFFSRPQX1MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFSRPQX0P5MA10TR (Q, D, CK, SN, R);
output Q;
input  D, CK, SN, R;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  not   XX1 (xRN, R);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$SN$Q  = 1.0,
    tphl$SN$Q  = 1.0,
    tplh$R$Q  = 1.0,
    tphl$R$Q  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tsetup$SN$CK    = 1.0,
    thold$SN$CK    = 0.5,
    tminpwl$SN     = 1.0,
    tminpwh$SN     = 1.0,
    tsetup$R$CK    = 1.0,
    thold$R$CK    = 0.5,
    tminpwl$R     = 1.0,
    tminpwh$R     = 1.0,
    thold$R$SN = 1.0,
    thold$SN$R = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK, negedge R &&& (SN == 1'b1), tsetup$R$CK, thold$R$CK, NOTIFIER);
    $width(posedge R &&& (SN == 1'b1), tminpwh$R, 0, NOTIFIER);
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK, thold$SN$CK, NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    $hold(negedge R, negedge SN, thold$SN$R, NOTIFIER);    
    $hold(posedge SN, posedge R, thold$R$SN, NOTIFIER);    
    if (D == 1'b0 && SN == 1'b1 && CK == 1'b0)
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b0 && R == 1'b0 && CK == 1'b0)
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q); 
    if (D == 1'b0 && SN == 1'b1 && CK == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b0 && R == 1'b0 && CK == 1'b1)
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q); 
    if (D == 1'b1 && SN == 1'b1 && CK == 1'b0)
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b1 && R == 1'b0 && CK == 1'b0)
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q); 
    if (D == 1'b1 && SN == 1'b1 && CK == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b1 && R == 1'b0 && CK == 1'b1)
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q); 

   endspecify
endmodule // DFFSRPQX0P5MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFSQNX3MA10TR (QN, D, CK, SN);
output QN;
input  D, CK, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$SN$QN  = 1.0,
    tphl$SN$QN  = 1.0,
    tplh$CK$QN	= 1.0,
    tphl$CK$QN	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    thold$SN$CK = 0.5,
    tsetup$SN$CK = 1.0,
    tminpwl$SN    = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (QN -: D)) = (tplh$CK$QN,   tphl$CK$QN);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK, thold$SN$CK, NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    if (D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b0)) = (tplh$SN$QN); 
    if (D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b0)) = (tplh$SN$QN); 
    if (D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b0)) = (tplh$SN$QN); 
    if (D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b0)) = (tplh$SN$QN); 

   endspecify
endmodule // DFFSQNX3MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFSQNX2MA10TR (QN, D, CK, SN);
output QN;
input  D, CK, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$SN$QN  = 1.0,
    tphl$SN$QN  = 1.0,
    tplh$CK$QN	= 1.0,
    tphl$CK$QN	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    thold$SN$CK = 0.5,
    tsetup$SN$CK = 1.0,
    tminpwl$SN    = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (QN -: D)) = (tplh$CK$QN,   tphl$CK$QN);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK, thold$SN$CK, NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    if (D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b0)) = (tplh$SN$QN); 
    if (D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b0)) = (tplh$SN$QN); 
    if (D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b0)) = (tplh$SN$QN); 
    if (D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b0)) = (tplh$SN$QN); 

   endspecify
endmodule // DFFSQNX2MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFSQNX1MA10TR (QN, D, CK, SN);
output QN;
input  D, CK, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$SN$QN  = 1.0,
    tphl$SN$QN  = 1.0,
    tplh$CK$QN	= 1.0,
    tphl$CK$QN	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    thold$SN$CK = 0.5,
    tsetup$SN$CK = 1.0,
    tminpwl$SN    = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (QN -: D)) = (tplh$CK$QN,   tphl$CK$QN);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK, thold$SN$CK, NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    if (D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b0)) = (tplh$SN$QN); 
    if (D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b0)) = (tplh$SN$QN); 
    if (D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b0)) = (tplh$SN$QN); 
    if (D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b0)) = (tplh$SN$QN); 

   endspecify
endmodule // DFFSQNX1MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFSQNX0P5MA10TR (QN, D, CK, SN);
output QN;
input  D, CK, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$SN$QN  = 1.0,
    tphl$SN$QN  = 1.0,
    tplh$CK$QN	= 1.0,
    tphl$CK$QN	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    thold$SN$CK = 0.5,
    tsetup$SN$CK = 1.0,
    tminpwl$SN    = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (QN -: D)) = (tplh$CK$QN,   tphl$CK$QN);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK, thold$SN$CK, NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    if (D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b0)) = (tplh$SN$QN); 
    if (D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b0)) = (tplh$SN$QN); 
    if (D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (QN -: 1'b0)) = (tplh$SN$QN); 
    if (D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (QN -: 1'b0)) = (tplh$SN$QN); 

   endspecify
endmodule // DFFSQNX0P5MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFSQX4MA10TR (Q, D, CK, SN);
output Q;
input  D, CK, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$SN$Q  = 1.0,
    tphl$SN$Q  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tsetup$SN$CK    = 1.0,
    thold$SN$CK    = 0.5,
    tminpwl$SN     = 1.0,
    tminpwh$SN     = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK, thold$SN$CK, NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    if (D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q);

   endspecify
endmodule // DFFSQX4MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFSQX3MA10TR (Q, D, CK, SN);
output Q;
input  D, CK, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$SN$Q  = 1.0,
    tphl$SN$Q  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tsetup$SN$CK    = 1.0,
    thold$SN$CK    = 0.5,
    tminpwl$SN     = 1.0,
    tminpwh$SN     = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK, thold$SN$CK, NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    if (D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q);

   endspecify
endmodule // DFFSQX3MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFSQX2MA10TR (Q, D, CK, SN);
output Q;
input  D, CK, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$SN$Q  = 1.0,
    tphl$SN$Q  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tsetup$SN$CK    = 1.0,
    thold$SN$CK    = 0.5,
    tminpwl$SN     = 1.0,
    tminpwh$SN     = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK, thold$SN$CK, NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    if (D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q);

   endspecify
endmodule // DFFSQX2MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFSQX1MA10TR (Q, D, CK, SN);
output Q;
input  D, CK, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$SN$Q  = 1.0,
    tphl$SN$Q  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tsetup$SN$CK    = 1.0,
    thold$SN$CK    = 0.5,
    tminpwl$SN     = 1.0,
    tminpwh$SN     = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK, thold$SN$CK, NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    if (D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q);

   endspecify
endmodule // DFFSQX1MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFSQX0P5MA10TR (Q, D, CK, SN);
output Q;
input  D, CK, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$SN$Q  = 1.0,
    tphl$SN$Q  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tsetup$SN$CK    = 1.0,
    thold$SN$CK    = 0.5,
    tminpwl$SN     = 1.0,
    tminpwh$SN     = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK, posedge SN, tsetup$SN$CK, thold$SN$CK, NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    if (D == 1'b0 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && CK == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b1 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q); 
    if (D == 1'b0 && CK == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q, tphl$SN$Q);

   endspecify
endmodule // DFFSQX0P5MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFRPQNX3MA10TR (QN, D, CK, R);
output QN;
input  D, CK, R;
reg NOTIFIER;
supply1 xSN;

  not   XX0 (xRN, R);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$R$QN  = 1.0,
    tphl$R$QN  = 1.0,
    tplh$CK$QN	= 1.0,
    tphl$CK$QN	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    thold$R$CK = 0.5,
    tsetup$R$CK = 1.0,
    tminpwh$R    = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (QN -: D)) = (tplh$CK$QN,   tphl$CK$QN);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK, negedge R, tsetup$R$CK, thold$R$CK, NOTIFIER);
    $width(posedge R, tminpwh$R, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    if (D == 1'b0 && CK == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = ( tphl$R$QN); 
    if (D == 1'b0 && CK == 1'b1 )
       (posedge  R *> (QN -: 1'b1)) = ( tphl$R$QN); 
    if (D == 1'b1 && CK == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = ( tphl$R$QN); 
    if (D == 1'b1 && CK == 1'b1 )
       (posedge  R *> (QN -: 1'b1)) = ( tphl$R$QN); 

   endspecify
endmodule // DFFRPQNX3MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFRPQNX2MA10TR (QN, D, CK, R);
output QN;
input  D, CK, R;
reg NOTIFIER;
supply1 xSN;

  not   XX0 (xRN, R);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$R$QN  = 1.0,
    tphl$R$QN  = 1.0,
    tplh$CK$QN	= 1.0,
    tphl$CK$QN	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    thold$R$CK = 0.5,
    tsetup$R$CK = 1.0,
    tminpwh$R    = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (QN -: D)) = (tplh$CK$QN,   tphl$CK$QN);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK, negedge R, tsetup$R$CK, thold$R$CK, NOTIFIER);
    $width(posedge R, tminpwh$R, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    if (D == 1'b0 && CK == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = ( tphl$R$QN); 
    if (D == 1'b0 && CK == 1'b1 )
       (posedge  R *> (QN -: 1'b1)) = ( tphl$R$QN); 
    if (D == 1'b1 && CK == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = ( tphl$R$QN); 
    if (D == 1'b1 && CK == 1'b1 )
       (posedge  R *> (QN -: 1'b1)) = ( tphl$R$QN); 

   endspecify
endmodule // DFFRPQNX2MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFRPQNX1MA10TR (QN, D, CK, R);
output QN;
input  D, CK, R;
reg NOTIFIER;
supply1 xSN;

  not   XX0 (xRN, R);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$R$QN  = 1.0,
    tphl$R$QN  = 1.0,
    tplh$CK$QN	= 1.0,
    tphl$CK$QN	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    thold$R$CK = 0.5,
    tsetup$R$CK = 1.0,
    tminpwh$R    = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (QN -: D)) = (tplh$CK$QN,   tphl$CK$QN);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK, negedge R, tsetup$R$CK, thold$R$CK, NOTIFIER);
    $width(posedge R, tminpwh$R, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    if (D == 1'b0 && CK == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = ( tphl$R$QN); 
    if (D == 1'b0 && CK == 1'b1 )
       (posedge  R *> (QN -: 1'b1)) = ( tphl$R$QN); 
    if (D == 1'b1 && CK == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = ( tphl$R$QN); 
    if (D == 1'b1 && CK == 1'b1 )
       (posedge  R *> (QN -: 1'b1)) = ( tphl$R$QN); 

   endspecify
endmodule // DFFRPQNX1MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFRPQNX0P5MA10TR (QN, D, CK, R);
output QN;
input  D, CK, R;
reg NOTIFIER;
supply1 xSN;

  not   XX0 (xRN, R);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$R$QN  = 1.0,
    tphl$R$QN  = 1.0,
    tplh$CK$QN	= 1.0,
    tphl$CK$QN	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    thold$R$CK = 0.5,
    tsetup$R$CK = 1.0,
    tminpwh$R    = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (QN -: D)) = (tplh$CK$QN,   tphl$CK$QN);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK, negedge R, tsetup$R$CK, thold$R$CK, NOTIFIER);
    $width(posedge R, tminpwh$R, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    if (D == 1'b0 && CK == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = ( tphl$R$QN); 
    if (D == 1'b0 && CK == 1'b1 )
       (posedge  R *> (QN -: 1'b1)) = ( tphl$R$QN); 
    if (D == 1'b1 && CK == 1'b0 )
       (posedge  R *> (QN -: 1'b1)) = ( tphl$R$QN); 
    if (D == 1'b1 && CK == 1'b1 )
       (posedge  R *> (QN -: 1'b1)) = ( tphl$R$QN); 

   endspecify
endmodule // DFFRPQNX0P5MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFRPQX4MA10TR (Q, D, CK, R);
output Q;
input  D, CK, R;
reg NOTIFIER;
supply1 xSN;

  not   XX0 (xRN, R);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$R$Q  = 1.0,
    tphl$R$Q  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tsetup$R$CK    = 1.0,
    thold$R$CK    = 0.5,
    tminpwl$R     = 1.0,
    tminpwh$R     = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK, negedge R, tsetup$R$CK, thold$R$CK, NOTIFIER);
    $width(posedge R, tminpwh$R, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    if (D == 1'b0 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b0 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b1 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b1 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 

   endspecify
endmodule // DFFRPQX4MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFRPQX3MA10TR (Q, D, CK, R);
output Q;
input  D, CK, R;
reg NOTIFIER;
supply1 xSN;

  not   XX0 (xRN, R);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$R$Q  = 1.0,
    tphl$R$Q  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tsetup$R$CK    = 1.0,
    thold$R$CK    = 0.5,
    tminpwl$R     = 1.0,
    tminpwh$R     = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK, negedge R, tsetup$R$CK, thold$R$CK, NOTIFIER);
    $width(posedge R, tminpwh$R, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    if (D == 1'b0 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b0 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b1 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b1 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 

   endspecify
endmodule // DFFRPQX3MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFRPQX2MA10TR (Q, D, CK, R);
output Q;
input  D, CK, R;
reg NOTIFIER;
supply1 xSN;

  not   XX0 (xRN, R);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$R$Q  = 1.0,
    tphl$R$Q  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tsetup$R$CK    = 1.0,
    thold$R$CK    = 0.5,
    tminpwl$R     = 1.0,
    tminpwh$R     = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK, negedge R, tsetup$R$CK, thold$R$CK, NOTIFIER);
    $width(posedge R, tminpwh$R, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    if (D == 1'b0 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b0 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b1 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b1 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 

   endspecify
endmodule // DFFRPQX2MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFRPQX1MA10TR (Q, D, CK, R);
output Q;
input  D, CK, R;
reg NOTIFIER;
supply1 xSN;

  not   XX0 (xRN, R);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$R$Q  = 1.0,
    tphl$R$Q  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tsetup$R$CK    = 1.0,
    thold$R$CK    = 0.5,
    tminpwl$R     = 1.0,
    tminpwh$R     = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK, negedge R, tsetup$R$CK, thold$R$CK, NOTIFIER);
    $width(posedge R, tminpwh$R, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    if (D == 1'b0 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b0 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b1 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b1 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 

   endspecify
endmodule // DFFRPQX1MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFRPQX0P5MA10TR (Q, D, CK, R);
output Q;
input  D, CK, R;
reg NOTIFIER;
supply1 xSN;

  not   XX0 (xRN, R);
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$R$Q  = 1.0,
    tphl$R$Q  = 1.0,
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tsetup$R$CK    = 1.0,
    thold$R$CK    = 0.5,
    tminpwl$R     = 1.0,
    tminpwh$R     = 1.0,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK, negedge R, tsetup$R$CK, thold$R$CK, NOTIFIER);
    $width(posedge R, tminpwh$R, 0, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);
    if (D == 1'b0 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b0 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b1 && CK == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b1 && CK == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 

   endspecify
endmodule // DFFRPQX0P5MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFQNX3MA10TR (QN, D, CK);
output QN;
input  D, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$CK$QN	= 1.0,
    tphl$CK$QN	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (QN -: D)) = (tplh$CK$QN,   tphl$CK$QN);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // DFFQNX3MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFQNX2MA10TR (QN, D, CK);
output QN;
input  D, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$CK$QN	= 1.0,
    tphl$CK$QN	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (QN -: D)) = (tplh$CK$QN,   tphl$CK$QN);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // DFFQNX2MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFQNX1MA10TR (QN, D, CK);
output QN;
input  D, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$CK$QN	= 1.0,
    tphl$CK$QN	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (QN -: D)) = (tplh$CK$QN,   tphl$CK$QN);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // DFFQNX1MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFQNX0P5MA10TR (QN, D, CK);
output QN;
input  D, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$CK$QN	= 1.0,
    tphl$CK$QN	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (QN -: D)) = (tplh$CK$QN,   tphl$CK$QN);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // DFFQNX0P5MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFQX4MA10TR (Q, D, CK);
output Q;
input  D, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // DFFQX4MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFQX3MA10TR (Q, D, CK);
output Q;
input  D, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // DFFQX3MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFQX2MA10TR (Q, D, CK);
output Q;
input  D, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // DFFQX2MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFQX1MA10TR (Q, D, CK);
output Q;
input  D, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // DFFQX1MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFQX0P5MA10TR (Q, D, CK);
output Q;
input  D, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$D$CK	= 1.0,
    thold$D$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;


    if (flag)
      (posedge CK *> (Q +: D)) = (tplh$CK$Q,    tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge D, tsetup$D$CK, thold$D$CK, NOTIFIER);
    $width(negedge CK &&& (flag == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag == 1), tminpwh$CK, 0, NOTIFIER); 
    $period(posedge CK &&& (flag == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // DFFQX0P5MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFNSRPQX3MA10TR (Q, D, CKN, SN, R);
output Q;
input  D, CKN, SN, R;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  not   XX1 (xRN, R);
  not     IC (clk, CKN);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$SN$Q  = 1.0,
    tphl$SN$Q  = 1.0,
    tplh$R$Q  = 1.0,
    tphl$R$Q  = 1.0,
    tplh$CKN$Q	= 1.0,
    tphl$CKN$Q	= 1.0,
    tsetup$D$CKN	= 1.0,
    thold$D$CKN	= 0.5,
    thold$SN$R = 0.5,
    thold$R$SN = 0.5,
    tsetup$SN$CKN    = 1.0,
    thold$SN$CKN    = 0.5,
    tminpwl$SN     = 1.0,
    tminpwh$SN     = 1.0,
    tsetup$R$CKN    = 1.0,
    thold$R$CKN    = 0.5,
    tminpwl$R     = 1.0,
    tminpwh$R     = 1.0,
    tminpwl$CKN    = 1.0,
    tminpwh$CKN    = 1.0,
    tperiod$CKN    = 1.0;

    if (flag)
      (negedge CKN *> (Q    +: D)) = (tplh$CKN$Q,    tphl$CKN$Q);
    $setuphold(negedge CKN &&& (flag == 1), posedge D, tsetup$D$CKN, thold$D$CKN, NOTIFIER);
    $setuphold(negedge CKN &&& (flag == 1), negedge D, tsetup$D$CKN, thold$D$CKN, NOTIFIER);
    $setuphold(negedge CKN, negedge R &&& (SN == 1'b1), tsetup$R$CKN, thold$R$CKN, NOTIFIER);
    $width(posedge R &&& (SN == 1'b1), tminpwh$R, 0, NOTIFIER);
    $setuphold(negedge CKN, posedge SN, tsetup$SN$CKN, thold$SN$CKN, NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $width(negedge CKN &&& (flag == 1), tminpwl$CKN, 0, NOTIFIER);
    $width(posedge CKN &&& (flag == 1), tminpwh$CKN, 0, NOTIFIER); 
    $period(posedge CKN &&& (flag == 1), tperiod$CKN, NOTIFIER);
    $hold(negedge R, negedge SN, thold$SN$R, NOTIFIER);    
    $hold(posedge SN, posedge R, thold$R$SN, NOTIFIER);    
    if (D == 1'b0 && SN == 1'b1 && CKN == 1'b0)
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b0 && R == 1'b0 && CKN == 1'b0)
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q); 
    if (D == 1'b0 && SN == 1'b1 && CKN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b0 && R == 1'b0 && CKN == 1'b1)
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q); 
    if (D == 1'b1 && SN == 1'b1 && CKN == 1'b0)
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b1 && R == 1'b0 && CKN == 1'b0)
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q); 
    if (D == 1'b1 && SN == 1'b1 && CKN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b1 && R == 1'b0 && CKN == 1'b1)
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q); 

   endspecify
endmodule // DFFNSRPQX3MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFNSRPQX2MA10TR (Q, D, CKN, SN, R);
output Q;
input  D, CKN, SN, R;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  not   XX1 (xRN, R);
  not     IC (clk, CKN);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$SN$Q  = 1.0,
    tphl$SN$Q  = 1.0,
    tplh$R$Q  = 1.0,
    tphl$R$Q  = 1.0,
    tplh$CKN$Q	= 1.0,
    tphl$CKN$Q	= 1.0,
    tsetup$D$CKN	= 1.0,
    thold$D$CKN	= 0.5,
    thold$SN$R = 0.5,
    thold$R$SN = 0.5,
    tsetup$SN$CKN    = 1.0,
    thold$SN$CKN    = 0.5,
    tminpwl$SN     = 1.0,
    tminpwh$SN     = 1.0,
    tsetup$R$CKN    = 1.0,
    thold$R$CKN    = 0.5,
    tminpwl$R     = 1.0,
    tminpwh$R     = 1.0,
    tminpwl$CKN    = 1.0,
    tminpwh$CKN    = 1.0,
    tperiod$CKN    = 1.0;

    if (flag)
      (negedge CKN *> (Q    +: D)) = (tplh$CKN$Q,    tphl$CKN$Q);
    $setuphold(negedge CKN &&& (flag == 1), posedge D, tsetup$D$CKN, thold$D$CKN, NOTIFIER);
    $setuphold(negedge CKN &&& (flag == 1), negedge D, tsetup$D$CKN, thold$D$CKN, NOTIFIER);
    $setuphold(negedge CKN, negedge R &&& (SN == 1'b1), tsetup$R$CKN, thold$R$CKN, NOTIFIER);
    $width(posedge R &&& (SN == 1'b1), tminpwh$R, 0, NOTIFIER);
    $setuphold(negedge CKN, posedge SN, tsetup$SN$CKN, thold$SN$CKN, NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $width(negedge CKN &&& (flag == 1), tminpwl$CKN, 0, NOTIFIER);
    $width(posedge CKN &&& (flag == 1), tminpwh$CKN, 0, NOTIFIER); 
    $period(posedge CKN &&& (flag == 1), tperiod$CKN, NOTIFIER);
    $hold(negedge R, negedge SN, thold$SN$R, NOTIFIER);    
    $hold(posedge SN, posedge R, thold$R$SN, NOTIFIER);    
    if (D == 1'b0 && SN == 1'b1 && CKN == 1'b0)
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b0 && R == 1'b0 && CKN == 1'b0)
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q); 
    if (D == 1'b0 && SN == 1'b1 && CKN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b0 && R == 1'b0 && CKN == 1'b1)
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q); 
    if (D == 1'b1 && SN == 1'b1 && CKN == 1'b0)
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b1 && R == 1'b0 && CKN == 1'b0)
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q); 
    if (D == 1'b1 && SN == 1'b1 && CKN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b1 && R == 1'b0 && CKN == 1'b1)
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q); 

   endspecify
endmodule // DFFNSRPQX2MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFNSRPQX1MA10TR (Q, D, CKN, SN, R);
output Q;
input  D, CKN, SN, R;
reg NOTIFIER;
  buf   XX0 (xSN, SN);
  not   XX1 (xRN, R);
  not     IC (clk, CKN);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$SN$Q  = 1.0,
    tphl$SN$Q  = 1.0,
    tplh$R$Q  = 1.0,
    tphl$R$Q  = 1.0,
    tplh$CKN$Q	= 1.0,
    tphl$CKN$Q	= 1.0,
    tsetup$D$CKN	= 1.0,
    thold$D$CKN	= 0.5,
    thold$SN$R = 0.5,
    thold$R$SN = 0.5,
    tsetup$SN$CKN    = 1.0,
    thold$SN$CKN    = 0.5,
    tminpwl$SN     = 1.0,
    tminpwh$SN     = 1.0,
    tsetup$R$CKN    = 1.0,
    thold$R$CKN    = 0.5,
    tminpwl$R     = 1.0,
    tminpwh$R     = 1.0,
    tminpwl$CKN    = 1.0,
    tminpwh$CKN    = 1.0,
    tperiod$CKN    = 1.0;

    if (flag)
      (negedge CKN *> (Q    +: D)) = (tplh$CKN$Q,    tphl$CKN$Q);
    $setuphold(negedge CKN &&& (flag == 1), posedge D, tsetup$D$CKN, thold$D$CKN, NOTIFIER);
    $setuphold(negedge CKN &&& (flag == 1), negedge D, tsetup$D$CKN, thold$D$CKN, NOTIFIER);
    $setuphold(negedge CKN, negedge R &&& (SN == 1'b1), tsetup$R$CKN, thold$R$CKN, NOTIFIER);
    $width(posedge R &&& (SN == 1'b1), tminpwh$R, 0, NOTIFIER);
    $setuphold(negedge CKN, posedge SN, tsetup$SN$CKN, thold$SN$CKN, NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $width(negedge CKN &&& (flag == 1), tminpwl$CKN, 0, NOTIFIER);
    $width(posedge CKN &&& (flag == 1), tminpwh$CKN, 0, NOTIFIER); 
    $period(posedge CKN &&& (flag == 1), tperiod$CKN, NOTIFIER);
    $hold(negedge R, negedge SN, thold$SN$R, NOTIFIER);    
    $hold(posedge SN, posedge R, thold$R$SN, NOTIFIER);    
    if (D == 1'b0 && SN == 1'b1 && CKN == 1'b0)
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b0 && R == 1'b0 && CKN == 1'b0)
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q); 
    if (D == 1'b0 && SN == 1'b1 && CKN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b0 && R == 1'b0 && CKN == 1'b1)
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q); 
    if (D == 1'b1 && SN == 1'b1 && CKN == 1'b0)
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b1 && R == 1'b0 && CKN == 1'b0)
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q); 
    if (D == 1'b1 && SN == 1'b1 && CKN == 1'b1)
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b1 && R == 1'b0 && CKN == 1'b1)
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q); 

   endspecify
endmodule // DFFNSRPQX1MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFNSQX3MA10TR (Q, D, CKN, SN);
output Q;
input  D, CKN, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  not     IC (clk, CKN);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$SN$Q  = 1.0,
    tphl$SN$Q  = 1.0,
    tplh$CKN$Q	= 1.0,
    tphl$CKN$Q	= 1.0,
    tsetup$D$CKN	= 1.0,
    thold$D$CKN	= 0.5,
    tsetup$SN$CKN    = 1.0,
    thold$SN$CKN    = 0.5,
    tminpwl$SN     = 1.0,
    tminpwh$SN     = 1.0,
    tminpwl$CKN    = 1.0,
    tminpwh$CKN    = 1.0,
    tperiod$CKN    = 1.0;

    if (flag)
      (negedge CKN *> (Q    +: D)) = (tplh$CKN$Q,    tphl$CKN$Q);
    $setuphold(negedge CKN &&& (flag == 1), posedge D, tsetup$D$CKN, thold$D$CKN, NOTIFIER);
    $setuphold(negedge CKN &&& (flag == 1), negedge D, tsetup$D$CKN, thold$D$CKN, NOTIFIER);
    $setuphold(negedge CKN, posedge SN, tsetup$SN$CKN, thold$SN$CKN, NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $width(negedge CKN &&& (flag == 1), tminpwl$CKN, 0, NOTIFIER);
    $width(posedge CKN &&& (flag == 1), tminpwh$CKN, 0, NOTIFIER); 
    $period(posedge CKN &&& (flag == 1), tperiod$CKN, NOTIFIER);
    if (D == 1'b0 && CKN == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q); 
    if (D == 1'b0 && CKN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q); 
    if (D == 1'b1 && CKN == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q); 
    if (D == 1'b1 && CKN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q); 

   endspecify
endmodule // DFFNSQX3MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFNSQX2MA10TR (Q, D, CKN, SN);
output Q;
input  D, CKN, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  not     IC (clk, CKN);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$SN$Q  = 1.0,
    tphl$SN$Q  = 1.0,
    tplh$CKN$Q	= 1.0,
    tphl$CKN$Q	= 1.0,
    tsetup$D$CKN	= 1.0,
    thold$D$CKN	= 0.5,
    tsetup$SN$CKN    = 1.0,
    thold$SN$CKN    = 0.5,
    tminpwl$SN     = 1.0,
    tminpwh$SN     = 1.0,
    tminpwl$CKN    = 1.0,
    tminpwh$CKN    = 1.0,
    tperiod$CKN    = 1.0;

    if (flag)
      (negedge CKN *> (Q    +: D)) = (tplh$CKN$Q,    tphl$CKN$Q);
    $setuphold(negedge CKN &&& (flag == 1), posedge D, tsetup$D$CKN, thold$D$CKN, NOTIFIER);
    $setuphold(negedge CKN &&& (flag == 1), negedge D, tsetup$D$CKN, thold$D$CKN, NOTIFIER);
    $setuphold(negedge CKN, posedge SN, tsetup$SN$CKN, thold$SN$CKN, NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $width(negedge CKN &&& (flag == 1), tminpwl$CKN, 0, NOTIFIER);
    $width(posedge CKN &&& (flag == 1), tminpwh$CKN, 0, NOTIFIER); 
    $period(posedge CKN &&& (flag == 1), tperiod$CKN, NOTIFIER);
    if (D == 1'b0 && CKN == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q); 
    if (D == 1'b0 && CKN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q); 
    if (D == 1'b1 && CKN == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q); 
    if (D == 1'b1 && CKN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q); 

   endspecify
endmodule // DFFNSQX2MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFNSQX1MA10TR (Q, D, CKN, SN);
output Q;
input  D, CKN, SN;
reg NOTIFIER;
supply1 xRN;

  buf   XX0 (xSN, SN);
  not     IC (clk, CKN);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$SN$Q  = 1.0,
    tphl$SN$Q  = 1.0,
    tplh$CKN$Q	= 1.0,
    tphl$CKN$Q	= 1.0,
    tsetup$D$CKN	= 1.0,
    thold$D$CKN	= 0.5,
    tsetup$SN$CKN    = 1.0,
    thold$SN$CKN    = 0.5,
    tminpwl$SN     = 1.0,
    tminpwh$SN     = 1.0,
    tminpwl$CKN    = 1.0,
    tminpwh$CKN    = 1.0,
    tperiod$CKN    = 1.0;

    if (flag)
      (negedge CKN *> (Q    +: D)) = (tplh$CKN$Q,    tphl$CKN$Q);
    $setuphold(negedge CKN &&& (flag == 1), posedge D, tsetup$D$CKN, thold$D$CKN, NOTIFIER);
    $setuphold(negedge CKN &&& (flag == 1), negedge D, tsetup$D$CKN, thold$D$CKN, NOTIFIER);
    $setuphold(negedge CKN, posedge SN, tsetup$SN$CKN, thold$SN$CKN, NOTIFIER);
    $width(negedge SN, tminpwl$SN, 0, NOTIFIER);
    $width(negedge CKN &&& (flag == 1), tminpwl$CKN, 0, NOTIFIER);
    $width(posedge CKN &&& (flag == 1), tminpwh$CKN, 0, NOTIFIER); 
    $period(posedge CKN &&& (flag == 1), tperiod$CKN, NOTIFIER);
    if (D == 1'b0 && CKN == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q); 
    if (D == 1'b0 && CKN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q); 
    if (D == 1'b1 && CKN == 1'b0 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q); 
    if (D == 1'b1 && CKN == 1'b1 )
       (negedge  SN *> (Q +: 1'b1)) = (tplh$SN$Q); 

   endspecify
endmodule // DFFNSQX1MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFNRPQX3MA10TR (Q, D, CKN, R);
output Q;
input  D, CKN, R;
reg NOTIFIER;
supply1 xSN;

  not   XX0 (xRN, R);
  not     IC (clk, CKN);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$R$Q  = 1.0,
    tphl$R$Q  = 1.0,
    tplh$CKN$Q	= 1.0,
    tphl$CKN$Q	= 1.0,
    tsetup$D$CKN	= 1.0,
    thold$D$CKN	= 0.5,
    tsetup$R$CKN    = 1.0,
    thold$R$CKN    = 0.5,
    tminpwl$R     = 1.0,
    tminpwh$R     = 1.0,
    tminpwl$CKN    = 1.0,
    tminpwh$CKN    = 1.0,
    tperiod$CKN    = 1.0;

    if (flag)
      (negedge CKN *> (Q    +: D)) = (tplh$CKN$Q,    tphl$CKN$Q);
    $setuphold(negedge CKN &&& (flag == 1), posedge D, tsetup$D$CKN, thold$D$CKN, NOTIFIER);
    $setuphold(negedge CKN &&& (flag == 1), negedge D, tsetup$D$CKN, thold$D$CKN, NOTIFIER);
    $setuphold(negedge CKN, negedge R , tsetup$R$CKN, thold$R$CKN, NOTIFIER);
    $width(posedge R , tminpwh$R, 0, NOTIFIER);
    $width(negedge CKN &&& (flag == 1), tminpwl$CKN, 0, NOTIFIER);
    $width(posedge CKN &&& (flag == 1), tminpwh$CKN, 0, NOTIFIER); 
    $period(posedge CKN &&& (flag == 1), tperiod$CKN, NOTIFIER);
    if (D == 1'b0 && CKN == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b0 && CKN == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b1 && CKN == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b1 && CKN == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 

   endspecify
endmodule // DFFNRPQX3MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFNRPQX2MA10TR (Q, D, CKN, R);
output Q;
input  D, CKN, R;
reg NOTIFIER;
supply1 xSN;

  not   XX0 (xRN, R);
  not     IC (clk, CKN);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$R$Q  = 1.0,
    tphl$R$Q  = 1.0,
    tplh$CKN$Q	= 1.0,
    tphl$CKN$Q	= 1.0,
    tsetup$D$CKN	= 1.0,
    thold$D$CKN	= 0.5,
    tsetup$R$CKN    = 1.0,
    thold$R$CKN    = 0.5,
    tminpwl$R     = 1.0,
    tminpwh$R     = 1.0,
    tminpwl$CKN    = 1.0,
    tminpwh$CKN    = 1.0,
    tperiod$CKN    = 1.0;

    if (flag)
      (negedge CKN *> (Q    +: D)) = (tplh$CKN$Q,    tphl$CKN$Q);
    $setuphold(negedge CKN &&& (flag == 1), posedge D, tsetup$D$CKN, thold$D$CKN, NOTIFIER);
    $setuphold(negedge CKN &&& (flag == 1), negedge D, tsetup$D$CKN, thold$D$CKN, NOTIFIER);
    $setuphold(negedge CKN, negedge R , tsetup$R$CKN, thold$R$CKN, NOTIFIER);
    $width(posedge R , tminpwh$R, 0, NOTIFIER);
    $width(negedge CKN &&& (flag == 1), tminpwl$CKN, 0, NOTIFIER);
    $width(posedge CKN &&& (flag == 1), tminpwh$CKN, 0, NOTIFIER); 
    $period(posedge CKN &&& (flag == 1), tperiod$CKN, NOTIFIER);
    if (D == 1'b0 && CKN == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b0 && CKN == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b1 && CKN == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b1 && CKN == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 

   endspecify
endmodule // DFFNRPQX2MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFNRPQX1MA10TR (Q, D, CKN, R);
output Q;
input  D, CKN, R;
reg NOTIFIER;
supply1 xSN;

  not   XX0 (xRN, R);
  not     IC (clk, CKN);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$R$Q  = 1.0,
    tphl$R$Q  = 1.0,
    tplh$CKN$Q	= 1.0,
    tphl$CKN$Q	= 1.0,
    tsetup$D$CKN	= 1.0,
    thold$D$CKN	= 0.5,
    tsetup$R$CKN    = 1.0,
    thold$R$CKN    = 0.5,
    tminpwl$R     = 1.0,
    tminpwh$R     = 1.0,
    tminpwl$CKN    = 1.0,
    tminpwh$CKN    = 1.0,
    tperiod$CKN    = 1.0;

    if (flag)
      (negedge CKN *> (Q    +: D)) = (tplh$CKN$Q,    tphl$CKN$Q);
    $setuphold(negedge CKN &&& (flag == 1), posedge D, tsetup$D$CKN, thold$D$CKN, NOTIFIER);
    $setuphold(negedge CKN &&& (flag == 1), negedge D, tsetup$D$CKN, thold$D$CKN, NOTIFIER);
    $setuphold(negedge CKN, negedge R , tsetup$R$CKN, thold$R$CKN, NOTIFIER);
    $width(posedge R , tminpwh$R, 0, NOTIFIER);
    $width(negedge CKN &&& (flag == 1), tminpwl$CKN, 0, NOTIFIER);
    $width(posedge CKN &&& (flag == 1), tminpwh$CKN, 0, NOTIFIER); 
    $period(posedge CKN &&& (flag == 1), tperiod$CKN, NOTIFIER);
    if (D == 1'b0 && CKN == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b0 && CKN == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b1 && CKN == 1'b0 )
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 
    if (D == 1'b1 && CKN == 1'b1 )
       (posedge  R *> (Q +: 1'b0)) = ( tphl$R$Q); 

   endspecify
endmodule // DFFNRPQX1MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFNQX3MA10TR (Q, D, CKN);
output Q;
input  D, CKN;
reg NOTIFIER;
supply1 xSN,xRN;
  not     IC (clk, CKN);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$CKN$Q	= 1.0,
    tphl$CKN$Q	= 1.0,
    tsetup$D$CKN	= 1.0,
    thold$D$CKN	= 0.5,
    tminpwl$CKN    = 1.0,
    tminpwh$CKN    = 1.0,
    tperiod$CKN    = 1.0;

    if (flag)
      (negedge CKN *> (Q    +: D)) = (tplh$CKN$Q,    tphl$CKN$Q);
    $setuphold(negedge CKN &&& (flag == 1), posedge D, tsetup$D$CKN, thold$D$CKN, NOTIFIER);
    $setuphold(negedge CKN &&& (flag == 1), negedge D, tsetup$D$CKN, thold$D$CKN, NOTIFIER);
    $width(negedge CKN &&& (flag == 1), tminpwl$CKN, 0, NOTIFIER);
    $width(posedge CKN &&& (flag == 1), tminpwh$CKN, 0, NOTIFIER); 
    $period(posedge CKN &&& (flag == 1), tperiod$CKN, NOTIFIER);

   endspecify
endmodule // DFFNQX3MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFNQX2MA10TR (Q, D, CKN);
output Q;
input  D, CKN;
reg NOTIFIER;
supply1 xSN,xRN;
  not     IC (clk, CKN);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$CKN$Q	= 1.0,
    tphl$CKN$Q	= 1.0,
    tsetup$D$CKN	= 1.0,
    thold$D$CKN	= 0.5,
    tminpwl$CKN    = 1.0,
    tminpwh$CKN    = 1.0,
    tperiod$CKN    = 1.0;

    if (flag)
      (negedge CKN *> (Q    +: D)) = (tplh$CKN$Q,    tphl$CKN$Q);
    $setuphold(negedge CKN &&& (flag == 1), posedge D, tsetup$D$CKN, thold$D$CKN, NOTIFIER);
    $setuphold(negedge CKN &&& (flag == 1), negedge D, tsetup$D$CKN, thold$D$CKN, NOTIFIER);
    $width(negedge CKN &&& (flag == 1), tminpwl$CKN, 0, NOTIFIER);
    $width(posedge CKN &&& (flag == 1), tminpwh$CKN, 0, NOTIFIER); 
    $period(posedge CKN &&& (flag == 1), tperiod$CKN, NOTIFIER);

   endspecify
endmodule // DFFNQX2MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module DFFNQX1MA10TR (Q, D, CKN);
output Q;
input  D, CKN;
reg NOTIFIER;
supply1 xSN,xRN;
  not     IC (clk, CKN);
  udp_dff I0 (n0, D, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$CKN$Q	= 1.0,
    tphl$CKN$Q	= 1.0,
    tsetup$D$CKN	= 1.0,
    thold$D$CKN	= 0.5,
    tminpwl$CKN    = 1.0,
    tminpwh$CKN    = 1.0,
    tperiod$CKN    = 1.0;

    if (flag)
      (negedge CKN *> (Q    +: D)) = (tplh$CKN$Q,    tphl$CKN$Q);
    $setuphold(negedge CKN &&& (flag == 1), posedge D, tsetup$D$CKN, thold$D$CKN, NOTIFIER);
    $setuphold(negedge CKN &&& (flag == 1), negedge D, tsetup$D$CKN, thold$D$CKN, NOTIFIER);
    $width(negedge CKN &&& (flag == 1), tminpwl$CKN, 0, NOTIFIER);
    $width(posedge CKN &&& (flag == 1), tminpwh$CKN, 0, NOTIFIER); 
    $period(posedge CKN &&& (flag == 1), tperiod$CKN, NOTIFIER);

   endspecify
endmodule // DFFNQX1MA10TR
`endcelldefine


//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFZX8MA10TR (Y, A, OE);
output Y;
input A, OE;

  bufif1 I0(Y, A, OE);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$OE$Y = 1.0,
      tphl$OE$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (OE *> Y) = (tplh$OE$Y, tphl$OE$Y);
  endspecify

endmodule // BUFZX8MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFZX6MA10TR (Y, A, OE);
output Y;
input A, OE;

  bufif1 I0(Y, A, OE);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$OE$Y = 1.0,
      tphl$OE$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (OE *> Y) = (tplh$OE$Y, tphl$OE$Y);
  endspecify

endmodule // BUFZX6MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFZX4MA10TR (Y, A, OE);
output Y;
input A, OE;

  bufif1 I0(Y, A, OE);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$OE$Y = 1.0,
      tphl$OE$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (OE *> Y) = (tplh$OE$Y, tphl$OE$Y);
  endspecify

endmodule // BUFZX4MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFZX3MA10TR (Y, A, OE);
output Y;
input A, OE;

  bufif1 I0(Y, A, OE);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$OE$Y = 1.0,
      tphl$OE$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (OE *> Y) = (tplh$OE$Y, tphl$OE$Y);
  endspecify

endmodule // BUFZX3MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFZX2MA10TR (Y, A, OE);
output Y;
input A, OE;

  bufif1 I0(Y, A, OE);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$OE$Y = 1.0,
      tphl$OE$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (OE *> Y) = (tplh$OE$Y, tphl$OE$Y);
  endspecify

endmodule // BUFZX2MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFZX1P4MA10TR (Y, A, OE);
output Y;
input A, OE;

  bufif1 I0(Y, A, OE);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$OE$Y = 1.0,
      tphl$OE$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (OE *> Y) = (tplh$OE$Y, tphl$OE$Y);
  endspecify

endmodule // BUFZX1P4MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFZX1MA10TR (Y, A, OE);
output Y;
input A, OE;

  bufif1 I0(Y, A, OE);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$OE$Y = 1.0,
      tphl$OE$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (OE *> Y) = (tplh$OE$Y, tphl$OE$Y);
  endspecify

endmodule // BUFZX1MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFZX16MA10TR (Y, A, OE);
output Y;
input A, OE;

  bufif1 I0(Y, A, OE);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$OE$Y = 1.0,
      tphl$OE$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (OE *> Y) = (tplh$OE$Y, tphl$OE$Y);
  endspecify

endmodule // BUFZX16MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFZX11MA10TR (Y, A, OE);
output Y;
input A, OE;

  bufif1 I0(Y, A, OE);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$OE$Y = 1.0,
      tphl$OE$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (OE *> Y) = (tplh$OE$Y, tphl$OE$Y);
  endspecify

endmodule // BUFZX11MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFHX9MA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFHX9MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFHX7P5MA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFHX7P5MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFHX6MA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFHX6MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFHX5MA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFHX5MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFHX4MA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFHX4MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFHX3P5MA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFHX3P5MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFHX3MA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFHX3MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFHX2P5MA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFHX2P5MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFHX2MA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFHX2MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFHX1P7MA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFHX1P7MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFHX1P4MA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFHX1P4MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFHX1P2MA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFHX1P2MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFHX1MA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFHX1MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFHX16MA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFHX16MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFHX13MA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFHX13MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFHX11MA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFHX11MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFHX0P8MA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFHX0P8MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFHX0P7MA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFHX0P7MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX9MA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX9MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX9BA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX9BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX7P5MA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX7P5MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX7P5BA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX7P5BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX6MA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX6MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX6BA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX6BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX5MA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX5MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX5BA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX5BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX4MA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX4MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX4BA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX4BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX3P5MA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX3P5MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX3P5BA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX3P5BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX3MA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX3MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX3BA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX3BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX2P5MA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX2P5MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX2P5BA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX2P5BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX2MA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX2MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX2BA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX2BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX1P7MA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX1P7MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX1P7BA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX1P7BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX1P4MA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX1P4MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX1P4BA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX1P4BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX1P2MA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX1P2MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX1P2BA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX1P2BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX1MA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX1MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX1BA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX1BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX16MA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX16MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX16BA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX16BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX13MA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX13MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX13BA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX13BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX11MA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX11MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX11BA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX11BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX0P8MA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX0P8MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX0P8BA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX0P8BA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX0P7MA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX0P7MA10TR
`endcelldefine
//$Id: buf.genpp,v 1.3 2006/01/20 11:16:19 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module BUFX0P7BA10TR (Y, A);
output Y;
input A;

  buf I0(Y, A);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
  endspecify

endmodule // BUFX0P7BA10TR
`endcelldefine
//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI32X6MA10TR (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;

  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$A2$Y = 1.0,
      tphl$A2$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // AOI32X6MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI32X4MA10TR (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;

  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$A2$Y = 1.0,
      tphl$A2$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // AOI32X4MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI32X3MA10TR (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;

  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$A2$Y = 1.0,
      tphl$A2$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // AOI32X3MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI32X2MA10TR (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;

  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$A2$Y = 1.0,
      tphl$A2$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // AOI32X2MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI32X1P4MA10TR (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;

  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$A2$Y = 1.0,
      tphl$A2$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // AOI32X1P4MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI32X1MA10TR (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;

  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$A2$Y = 1.0,
      tphl$A2$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // AOI32X1MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI32X0P7MA10TR (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;

  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$A2$Y = 1.0,
      tphl$A2$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // AOI32X0P7MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI32X0P5MA10TR (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;

  and I0(outA, A0, A1, A2);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$A2$Y = 1.0,
      tphl$A2$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && A2 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (A1 == 1'b1 && A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // AOI32X0P5MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI31X6MA10TR (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;

  and I0(outA, A0, A1, A2);
  nor I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$A2$Y = 1.0,
      tphl$A2$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
      (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y);
    if (A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AOI31X6MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI31X4MA10TR (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;

  and I0(outA, A0, A1, A2);
  nor I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$A2$Y = 1.0,
      tphl$A2$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
      (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y);
    if (A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AOI31X4MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI31X3MA10TR (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;

  and I0(outA, A0, A1, A2);
  nor I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$A2$Y = 1.0,
      tphl$A2$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
      (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y);
    if (A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AOI31X3MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI31X2MA10TR (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;

  and I0(outA, A0, A1, A2);
  nor I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$A2$Y = 1.0,
      tphl$A2$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
      (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y);
    if (A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AOI31X2MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI31X1P4MA10TR (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;

  and I0(outA, A0, A1, A2);
  nor I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$A2$Y = 1.0,
      tphl$A2$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
      (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y);
    if (A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AOI31X1P4MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI31X1MA10TR (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;

  and I0(outA, A0, A1, A2);
  nor I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$A2$Y = 1.0,
      tphl$A2$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
      (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y);
    if (A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AOI31X1MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI31X0P7MA10TR (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;

  and I0(outA, A0, A1, A2);
  nor I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$A2$Y = 1.0,
      tphl$A2$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
      (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y);
    if (A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AOI31X0P7MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI31X0P5MA10TR (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;

  and I0(outA, A0, A1, A2);
  nor I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$A2$Y = 1.0,
      tphl$A2$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
      (A2 *> Y) = (tplh$A2$Y, tphl$A2$Y);
    if (A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && A2 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AOI31X0P5MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI2XB1X8MA10TR (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;

  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor I2(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);
    if (A0 == 1'b1 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AOI2XB1X8MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI2XB1X6MA10TR (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;

  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor I2(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);
    if (A0 == 1'b1 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AOI2XB1X6MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI2XB1X4MA10TR (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;

  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor I2(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);
    if (A0 == 1'b1 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AOI2XB1X4MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI2XB1X3MA10TR (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;

  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor I2(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);
    if (A0 == 1'b1 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AOI2XB1X3MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI2XB1X2MA10TR (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;

  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor I2(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);
    if (A0 == 1'b1 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AOI2XB1X2MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI2XB1X1P4MA10TR (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;

  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor I2(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);
    if (A0 == 1'b1 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AOI2XB1X1P4MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI2XB1X1MA10TR (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;

  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor I2(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);
    if (A0 == 1'b1 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AOI2XB1X1MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI2XB1X0P7MA10TR (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;

  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor I2(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);
    if (A0 == 1'b1 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AOI2XB1X0P7MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI2XB1X0P5MA10TR (Y, A0, A1N, B0);
output Y;
input A0, A1N, B0;

  not I0 (outA1, A1N);
  and I1 (outA, A0, outA1);
  nor I2(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1N$Y = 1.0,
      tphl$A1N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1N *> Y) = (tplh$A1N$Y, tphl$A1N$Y);
    if (A0 == 1'b1 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1N == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1N == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AOI2XB1X0P5MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI22X8MA10TR (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // AOI22X8MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI22X6MA10TR (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // AOI22X6MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI22X4MA10TR (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // AOI22X4MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI22X3MA10TR (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // AOI22X3MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI22X2MA10TR (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // AOI22X2MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI22X1P4MA10TR (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // AOI22X1P4MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI22X1MA10TR (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // AOI22X1MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI22X0P7MA10TR (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // AOI22X0P7MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI22X0P5MA10TR (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // AOI22X0P5MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI222X4MA10TR (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;

  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor I3(Y, outA, outB, outC);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0,
      tplh$C1$Y = 1.0,
      tphl$C1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y);

  endspecify
endmodule // AOI222X4MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI222X3MA10TR (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;

  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor I3(Y, outA, outB, outC);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0,
      tplh$C1$Y = 1.0,
      tphl$C1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y);

  endspecify
endmodule // AOI222X3MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI222X2MA10TR (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;

  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor I3(Y, outA, outB, outC);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0,
      tplh$C1$Y = 1.0,
      tphl$C1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y);

  endspecify
endmodule // AOI222X2MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI222X1P4MA10TR (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;

  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor I3(Y, outA, outB, outC);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0,
      tplh$C1$Y = 1.0,
      tphl$C1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y);

  endspecify
endmodule // AOI222X1P4MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI222X1MA10TR (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;

  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor I3(Y, outA, outB, outC);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0,
      tplh$C1$Y = 1.0,
      tphl$C1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y);

  endspecify
endmodule // AOI222X1MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI222X0P7MA10TR (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;

  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor I3(Y, outA, outB, outC);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0,
      tplh$C1$Y = 1.0,
      tphl$C1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y);

  endspecify
endmodule // AOI222X0P7MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI222X0P5MA10TR (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;

  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  and I2(outC, C0, C1);
  nor I3(Y, outA, outB, outC);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0,
      tplh$C1$Y = 1.0,
      tphl$C1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 && C1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b1 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 && C1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b1 )
       (C1 *> Y) = (tplh$C1$Y, tphl$C1$Y);

  endspecify
endmodule // AOI222X0P5MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI221X4MA10TR (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;

  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, C0, outB, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && C0 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // AOI221X4MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI221X3MA10TR (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;

  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, C0, outB, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && C0 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // AOI221X3MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI221X2MA10TR (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;

  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, C0, outB, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && C0 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // AOI221X2MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI221X1P4MA10TR (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;

  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, C0, outB, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && C0 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // AOI221X1P4MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI221X1MA10TR (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;

  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, C0, outB, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && C0 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // AOI221X1MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI221X0P7MA10TR (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;

  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, C0, outB, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && C0 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // AOI221X0P7MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI221X0P5MA10TR (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;

  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  nor I2(Y, C0, outB, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 && C0 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 && C0 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B1 == 1'b1 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B1 == 1'b1 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && C0 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && C0 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b1 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 && B1 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // AOI221X0P5MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI21BX8MA10TR (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;

  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor I3 (Y,outA,outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0N$Y = 1.0,
      tphl$B0N$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y);

  endspecify
endmodule // AOI21BX8MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI21BX6MA10TR (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;

  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor I3 (Y,outA,outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0N$Y = 1.0,
      tphl$B0N$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y);

  endspecify
endmodule // AOI21BX6MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI21BX4MA10TR (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;

  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor I3 (Y,outA,outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0N$Y = 1.0,
      tphl$B0N$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y);

  endspecify
endmodule // AOI21BX4MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI21BX3MA10TR (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;

  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor I3 (Y,outA,outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0N$Y = 1.0,
      tphl$B0N$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y);

  endspecify
endmodule // AOI21BX3MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI21BX2MA10TR (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;

  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor I3 (Y,outA,outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0N$Y = 1.0,
      tphl$B0N$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y);

  endspecify
endmodule // AOI21BX2MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI21BX1P4MA10TR (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;

  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor I3 (Y,outA,outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0N$Y = 1.0,
      tphl$B0N$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y);

  endspecify
endmodule // AOI21BX1P4MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI21BX1MA10TR (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;

  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor I3 (Y,outA,outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0N$Y = 1.0,
      tphl$B0N$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y);

  endspecify
endmodule // AOI21BX1MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI21BX0P7MA10TR (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;

  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor I3 (Y,outA,outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0N$Y = 1.0,
      tphl$B0N$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y);

  endspecify
endmodule // AOI21BX0P7MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI21BX0P5MA10TR (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;

  and I0(outA, A0, A1);
  not I1 (outB, B0N);
  nor I3 (Y,outA,outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0N$Y = 1.0,
      tphl$B0N$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 )
       (B0N *> Y) = (tplh$B0N$Y, tphl$B0N$Y);

  endspecify
endmodule // AOI21BX0P5MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI21X8MA10TR (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  and I0(outA, A0, A1);
  nor I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AOI21X8MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI21X6MA10TR (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  and I0(outA, A0, A1);
  nor I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AOI21X6MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI21X4MA10TR (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  and I0(outA, A0, A1);
  nor I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AOI21X4MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI21X3MA10TR (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  and I0(outA, A0, A1);
  nor I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AOI21X3MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI21X2MA10TR (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  and I0(outA, A0, A1);
  nor I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AOI21X2MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI21X1P4MA10TR (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  and I0(outA, A0, A1);
  nor I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AOI21X1P4MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI21X1MA10TR (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  and I0(outA, A0, A1);
  nor I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AOI21X1MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI21X0P7MA10TR (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  and I0(outA, A0, A1);
  nor I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AOI21X0P7MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI21X0P5MA10TR (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  and I0(outA, A0, A1);
  nor I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AOI21X0P5MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI211X4MA10TR (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;

  and I0(outA, A0, A1);
  nor I1(Y, B0, C0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b0 && A1 == 1'b0 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // AOI211X4MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI211X3MA10TR (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;

  and I0(outA, A0, A1);
  nor I1(Y, B0, C0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b0 && A1 == 1'b0 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // AOI211X3MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI211X2MA10TR (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;

  and I0(outA, A0, A1);
  nor I1(Y, B0, C0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b0 && A1 == 1'b0 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // AOI211X2MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI211X1P4MA10TR (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;

  and I0(outA, A0, A1);
  nor I1(Y, B0, C0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b0 && A1 == 1'b0 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // AOI211X1P4MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI211X1MA10TR (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;

  and I0(outA, A0, A1);
  nor I1(Y, B0, C0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b0 && A1 == 1'b0 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // AOI211X1MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI211X0P7MA10TR (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;

  and I0(outA, A0, A1);
  nor I1(Y, B0, C0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b0 && A1 == 1'b0 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // AOI211X0P7MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AOI211X0P5MA10TR (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;

  and I0(outA, A0, A1);
  nor I1(Y, B0, C0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$C0$Y = 1.0,
      tphl$C0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b0 && A1 == 1'b0 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && C0 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 && B0 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 && B0 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y); 
    if (A0 == 1'b1 && A1 == 1'b0 && B0 == 1'b0 )
       (C0 *> Y) = (tplh$C0$Y, tphl$C0$Y);

  endspecify
endmodule // AOI211X0P5MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO22X6MA10TR (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  or I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // AO22X6MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO22X4MA10TR (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  or I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // AO22X4MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO22X3MA10TR (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  or I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // AO22X3MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO22X2MA10TR (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  or I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // AO22X2MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO22X1P4MA10TR (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  or I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // AO22X1P4MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO22X1MA10TR (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  or I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // AO22X1MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO22X0P7MA10TR (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  or I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // AO22X0P7MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO22X0P5MA10TR (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;

  and I0(outA, A0, A1);
  and I1(outB, B0, B1);
  or I2(Y, outA, outB);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
    if (A1 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A1 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y); 
    if (A0 == 1'b1 && B0 == 1'b1 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b1 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (A0 == 1'b1 && B0 == 1'b0 && B1 == 1'b0 )
       (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y); 
    if (B1 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B1 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (B0 == 1'b1 && A0 == 1'b1 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b1 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y); 
    if (B0 == 1'b1 && A0 == 1'b0 && A1 == 1'b0 )
       (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

  endspecify
endmodule // AO22X0P5MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO21BX6MA10TR (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;

  and I0(outA, A0, A1);
  not I1(outB, B0N);
  or I2(Y, outB, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0N$Y = 1.0,
      tphl$B0N$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
   if ( A0 == 1'b1 && A1 == 1'b0  )
      ( B0N *> Y) = ( tplh$B0N$Y, tphl$B0N$Y);
   if ( A0 == 1'b0 && A1 == 1'b1  )
      ( B0N *> Y) = ( tplh$B0N$Y, tphl$B0N$Y);
   if ( A0 == 1'b0 && A1 == 1'b0  )
      ( B0N *> Y) = ( tplh$B0N$Y, tphl$B0N$Y);

  endspecify
endmodule // AO21BX6MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO21BX4MA10TR (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;

  and I0(outA, A0, A1);
  not I1(outB, B0N);
  or I2(Y, outB, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0N$Y = 1.0,
      tphl$B0N$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
   if ( A0 == 1'b1 && A1 == 1'b0  )
      ( B0N *> Y) = ( tplh$B0N$Y, tphl$B0N$Y);
   if ( A0 == 1'b0 && A1 == 1'b1  )
      ( B0N *> Y) = ( tplh$B0N$Y, tphl$B0N$Y);
   if ( A0 == 1'b0 && A1 == 1'b0  )
      ( B0N *> Y) = ( tplh$B0N$Y, tphl$B0N$Y);

  endspecify
endmodule // AO21BX4MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO21BX3MA10TR (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;

  and I0(outA, A0, A1);
  not I1(outB, B0N);
  or I2(Y, outB, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0N$Y = 1.0,
      tphl$B0N$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
   if ( A0 == 1'b1 && A1 == 1'b0  )
      ( B0N *> Y) = ( tplh$B0N$Y, tphl$B0N$Y);
   if ( A0 == 1'b0 && A1 == 1'b1  )
      ( B0N *> Y) = ( tplh$B0N$Y, tphl$B0N$Y);
   if ( A0 == 1'b0 && A1 == 1'b0  )
      ( B0N *> Y) = ( tplh$B0N$Y, tphl$B0N$Y);

  endspecify
endmodule // AO21BX3MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO21BX2MA10TR (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;

  and I0(outA, A0, A1);
  not I1(outB, B0N);
  or I2(Y, outB, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0N$Y = 1.0,
      tphl$B0N$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
   if ( A0 == 1'b1 && A1 == 1'b0  )
      ( B0N *> Y) = ( tplh$B0N$Y, tphl$B0N$Y);
   if ( A0 == 1'b0 && A1 == 1'b1  )
      ( B0N *> Y) = ( tplh$B0N$Y, tphl$B0N$Y);
   if ( A0 == 1'b0 && A1 == 1'b0  )
      ( B0N *> Y) = ( tplh$B0N$Y, tphl$B0N$Y);

  endspecify
endmodule // AO21BX2MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO21BX1P4MA10TR (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;

  and I0(outA, A0, A1);
  not I1(outB, B0N);
  or I2(Y, outB, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0N$Y = 1.0,
      tphl$B0N$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
   if ( A0 == 1'b1 && A1 == 1'b0  )
      ( B0N *> Y) = ( tplh$B0N$Y, tphl$B0N$Y);
   if ( A0 == 1'b0 && A1 == 1'b1  )
      ( B0N *> Y) = ( tplh$B0N$Y, tphl$B0N$Y);
   if ( A0 == 1'b0 && A1 == 1'b0  )
      ( B0N *> Y) = ( tplh$B0N$Y, tphl$B0N$Y);

  endspecify
endmodule // AO21BX1P4MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO21BX1MA10TR (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;

  and I0(outA, A0, A1);
  not I1(outB, B0N);
  or I2(Y, outB, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0N$Y = 1.0,
      tphl$B0N$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
   if ( A0 == 1'b1 && A1 == 1'b0  )
      ( B0N *> Y) = ( tplh$B0N$Y, tphl$B0N$Y);
   if ( A0 == 1'b0 && A1 == 1'b1  )
      ( B0N *> Y) = ( tplh$B0N$Y, tphl$B0N$Y);
   if ( A0 == 1'b0 && A1 == 1'b0  )
      ( B0N *> Y) = ( tplh$B0N$Y, tphl$B0N$Y);

  endspecify
endmodule // AO21BX1MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO21BX0P7MA10TR (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;

  and I0(outA, A0, A1);
  not I1(outB, B0N);
  or I2(Y, outB, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0N$Y = 1.0,
      tphl$B0N$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
   if ( A0 == 1'b1 && A1 == 1'b0  )
      ( B0N *> Y) = ( tplh$B0N$Y, tphl$B0N$Y);
   if ( A0 == 1'b0 && A1 == 1'b1  )
      ( B0N *> Y) = ( tplh$B0N$Y, tphl$B0N$Y);
   if ( A0 == 1'b0 && A1 == 1'b0  )
      ( B0N *> Y) = ( tplh$B0N$Y, tphl$B0N$Y);

  endspecify
endmodule // AO21BX0P7MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO21BX0P5MA10TR (Y, A0, A1, B0N);
output Y;
input A0, A1, B0N;

  and I0(outA, A0, A1);
  not I1(outB, B0N);
  or I2(Y, outB, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0N$Y = 1.0,
      tphl$B0N$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
   if ( A0 == 1'b1 && A1 == 1'b0  )
      ( B0N *> Y) = ( tplh$B0N$Y, tphl$B0N$Y);
   if ( A0 == 1'b0 && A1 == 1'b1  )
      ( B0N *> Y) = ( tplh$B0N$Y, tphl$B0N$Y);
   if ( A0 == 1'b0 && A1 == 1'b0  )
      ( B0N *> Y) = ( tplh$B0N$Y, tphl$B0N$Y);

  endspecify
endmodule // AO21BX0P5MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO21X6MA10TR (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  and I0(outA, A0, A1);
  or I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AO21X6MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO21X4MA10TR (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  and I0(outA, A0, A1);
  or I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AO21X4MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO21X3MA10TR (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  and I0(outA, A0, A1);
  or I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AO21X3MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO21X2MA10TR (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  and I0(outA, A0, A1);
  or I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AO21X2MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO21X1P4MA10TR (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  and I0(outA, A0, A1);
  or I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AO21X1P4MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO21X1MA10TR (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  and I0(outA, A0, A1);
  or I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AO21X1MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO21X0P7MA10TR (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  and I0(outA, A0, A1);
  or I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AO21X0P7MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO21X0P5MA10TR (Y, A0, A1, B0);
output Y;
input A0, A1, B0;

  and I0(outA, A0, A1);
  or I1(Y, B0, outA);
  specify
    // delay parameters
    specparam
      tplh$A0$Y = 1.0,
      tphl$A0$Y = 1.0,
      tplh$A1$Y = 1.0,
      tphl$A1$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0;

    // path delays
      (A0 *> Y) = (tplh$A0$Y, tphl$A0$Y);
      (A1 *> Y) = (tplh$A1$Y, tphl$A1$Y);
    if (A0 == 1'b1 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b1 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y); 
    if (A0 == 1'b0 && A1 == 1'b0 )
       (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);

  endspecify
endmodule // AO21X0P5MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO1B2X6MA10TR (Y, A0N, B0, B1);
output Y;
input A0N, B0, B1;

  nand I1 (outB, B0, B1);
  nand I2 (Y, A0N, outB);
  specify
    // delay parameters
    specparam
      tplh$A0N$Y = 1.0,
      tphl$A0N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
      (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);
      (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

    if ( B0==1'b0 && B1==1'b0  ) 
       ( A0N *> Y ) = ( tplh$A0N$Y,  tphl$A0N$Y);
    if ( B0==1'b0 && B1==1'b1  ) 
       ( A0N *> Y ) = ( tplh$A0N$Y,  tphl$A0N$Y);
    if ( B0==1'b1 && B1==1'b0  ) 
       ( A0N *> Y ) = ( tplh$A0N$Y,  tphl$A0N$Y);
  endspecify
endmodule // AO1B2X6MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO1B2X4MA10TR (Y, A0N, B0, B1);
output Y;
input A0N, B0, B1;

  nand I1 (outB, B0, B1);
  nand I2 (Y, A0N, outB);
  specify
    // delay parameters
    specparam
      tplh$A0N$Y = 1.0,
      tphl$A0N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
      (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);
      (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

    if ( B0==1'b0 && B1==1'b0  ) 
       ( A0N *> Y ) = ( tplh$A0N$Y,  tphl$A0N$Y);
    if ( B0==1'b0 && B1==1'b1  ) 
       ( A0N *> Y ) = ( tplh$A0N$Y,  tphl$A0N$Y);
    if ( B0==1'b1 && B1==1'b0  ) 
       ( A0N *> Y ) = ( tplh$A0N$Y,  tphl$A0N$Y);
  endspecify
endmodule // AO1B2X4MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO1B2X3MA10TR (Y, A0N, B0, B1);
output Y;
input A0N, B0, B1;

  nand I1 (outB, B0, B1);
  nand I2 (Y, A0N, outB);
  specify
    // delay parameters
    specparam
      tplh$A0N$Y = 1.0,
      tphl$A0N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
      (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);
      (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

    if ( B0==1'b0 && B1==1'b0  ) 
       ( A0N *> Y ) = ( tplh$A0N$Y,  tphl$A0N$Y);
    if ( B0==1'b0 && B1==1'b1  ) 
       ( A0N *> Y ) = ( tplh$A0N$Y,  tphl$A0N$Y);
    if ( B0==1'b1 && B1==1'b0  ) 
       ( A0N *> Y ) = ( tplh$A0N$Y,  tphl$A0N$Y);
  endspecify
endmodule // AO1B2X3MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO1B2X2MA10TR (Y, A0N, B0, B1);
output Y;
input A0N, B0, B1;

  nand I1 (outB, B0, B1);
  nand I2 (Y, A0N, outB);
  specify
    // delay parameters
    specparam
      tplh$A0N$Y = 1.0,
      tphl$A0N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
      (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);
      (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

    if ( B0==1'b0 && B1==1'b0  ) 
       ( A0N *> Y ) = ( tplh$A0N$Y,  tphl$A0N$Y);
    if ( B0==1'b0 && B1==1'b1  ) 
       ( A0N *> Y ) = ( tplh$A0N$Y,  tphl$A0N$Y);
    if ( B0==1'b1 && B1==1'b0  ) 
       ( A0N *> Y ) = ( tplh$A0N$Y,  tphl$A0N$Y);
  endspecify
endmodule // AO1B2X2MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO1B2X1P4MA10TR (Y, A0N, B0, B1);
output Y;
input A0N, B0, B1;

  nand I1 (outB, B0, B1);
  nand I2 (Y, A0N, outB);
  specify
    // delay parameters
    specparam
      tplh$A0N$Y = 1.0,
      tphl$A0N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
      (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);
      (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

    if ( B0==1'b0 && B1==1'b0  ) 
       ( A0N *> Y ) = ( tplh$A0N$Y,  tphl$A0N$Y);
    if ( B0==1'b0 && B1==1'b1  ) 
       ( A0N *> Y ) = ( tplh$A0N$Y,  tphl$A0N$Y);
    if ( B0==1'b1 && B1==1'b0  ) 
       ( A0N *> Y ) = ( tplh$A0N$Y,  tphl$A0N$Y);
  endspecify
endmodule // AO1B2X1P4MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO1B2X1MA10TR (Y, A0N, B0, B1);
output Y;
input A0N, B0, B1;

  nand I1 (outB, B0, B1);
  nand I2 (Y, A0N, outB);
  specify
    // delay parameters
    specparam
      tplh$A0N$Y = 1.0,
      tphl$A0N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
      (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);
      (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

    if ( B0==1'b0 && B1==1'b0  ) 
       ( A0N *> Y ) = ( tplh$A0N$Y,  tphl$A0N$Y);
    if ( B0==1'b0 && B1==1'b1  ) 
       ( A0N *> Y ) = ( tplh$A0N$Y,  tphl$A0N$Y);
    if ( B0==1'b1 && B1==1'b0  ) 
       ( A0N *> Y ) = ( tplh$A0N$Y,  tphl$A0N$Y);
  endspecify
endmodule // AO1B2X1MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO1B2X0P7MA10TR (Y, A0N, B0, B1);
output Y;
input A0N, B0, B1;

  nand I1 (outB, B0, B1);
  nand I2 (Y, A0N, outB);
  specify
    // delay parameters
    specparam
      tplh$A0N$Y = 1.0,
      tphl$A0N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
      (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);
      (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

    if ( B0==1'b0 && B1==1'b0  ) 
       ( A0N *> Y ) = ( tplh$A0N$Y,  tphl$A0N$Y);
    if ( B0==1'b0 && B1==1'b1  ) 
       ( A0N *> Y ) = ( tplh$A0N$Y,  tphl$A0N$Y);
    if ( B0==1'b1 && B1==1'b0  ) 
       ( A0N *> Y ) = ( tplh$A0N$Y,  tphl$A0N$Y);
  endspecify
endmodule // AO1B2X0P7MA10TR
`endcelldefine





//$Id: aoi.genpp,v 1.9 2006/06/13 06:07:04 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AO1B2X0P5MA10TR (Y, A0N, B0, B1);
output Y;
input A0N, B0, B1;

  nand I1 (outB, B0, B1);
  nand I2 (Y, A0N, outB);
  specify
    // delay parameters
    specparam
      tplh$A0N$Y = 1.0,
      tphl$A0N$Y = 1.0,
      tplh$B0$Y = 1.0,
      tphl$B0$Y = 1.0,
      tplh$B1$Y = 1.0,
      tphl$B1$Y = 1.0;

    // path delays
      (B0 *> Y) = (tplh$B0$Y, tphl$B0$Y);
      (B1 *> Y) = (tplh$B1$Y, tphl$B1$Y);

    if ( B0==1'b0 && B1==1'b0  ) 
       ( A0N *> Y ) = ( tplh$A0N$Y,  tphl$A0N$Y);
    if ( B0==1'b0 && B1==1'b1  ) 
       ( A0N *> Y ) = ( tplh$A0N$Y,  tphl$A0N$Y);
    if ( B0==1'b1 && B1==1'b0  ) 
       ( A0N *> Y ) = ( tplh$A0N$Y,  tphl$A0N$Y);
  endspecify
endmodule // AO1B2X0P5MA10TR
`endcelldefine





//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AND4X8MA10TR (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // AND4X8MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AND4X6MA10TR (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // AND4X6MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AND4X4MA10TR (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // AND4X4MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AND4X3MA10TR (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // AND4X3MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AND4X2MA10TR (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // AND4X2MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AND4X1P4MA10TR (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // AND4X1P4MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AND4X1MA10TR (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // AND4X1MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AND4X0P7MA10TR (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // AND4X0P7MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AND4X0P5MA10TR (Y, A, B, C, D);
output Y;
input A, B, C, D;

  and (Y, A, B, C, D);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0,
      tplh$D$Y = 1.0,
      tphl$D$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
    (D *> Y) = (tplh$D$Y, tphl$D$Y);
  endspecify
endmodule // AND4X0P5MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AND3X8MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  and (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // AND3X8MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AND3X6MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  and (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // AND3X6MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AND3X4MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  and (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // AND3X4MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AND3X3MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  and (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // AND3X3MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AND3X2MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  and (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // AND3X2MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AND3X1P4MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  and (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // AND3X1P4MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AND3X1MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  and (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // AND3X1MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AND3X11MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  and (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // AND3X11MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AND3X0P7MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  and (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // AND3X0P7MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AND3X0P5MA10TR (Y, A, B, C);
output Y;
input A, B, C;

  and (Y, A, B, C);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0,
      tplh$C$Y = 1.0,
      tphl$C$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
    (C *> Y) = (tplh$C$Y, tphl$C$Y);
  endspecify
endmodule // AND3X0P5MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AND2X8MA10TR (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // AND2X8MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AND2X6MA10TR (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // AND2X6MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AND2X4MA10TR (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // AND2X4MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AND2X3MA10TR (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // AND2X3MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AND2X2MA10TR (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // AND2X2MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AND2X1P4MA10TR (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // AND2X1P4MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AND2X1MA10TR (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // AND2X1MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AND2X11MA10TR (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // AND2X11MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AND2X0P7MA10TR (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // AND2X0P7MA10TR
`endcelldefine
//$Id: comb.genpp,v 1.5 2006/06/13 06:01:59 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module AND2X0P5MA10TR (Y, A, B);
output Y;
input A, B;

  and (Y, A, B);
  specify
    // delay parameters
    specparam
      tplh$A$Y = 1.0,
      tphl$A$Y = 1.0,
      tplh$B$Y = 1.0,
      tphl$B$Y = 1.0;

    // path delays
    (A *> Y) = (tplh$A$Y, tphl$A$Y);
    (B *> Y) = (tplh$B$Y, tphl$B$Y);
  endspecify
endmodule // AND2X0P5MA10TR
`endcelldefine
//$Id: add.genpp,v 1.7 2006/06/01 15:56:41 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module ADDHX2MA10TR ( S, CO, A, B);
output S, CO;
input A, B;
  xor I0(S, A, B);
  and I1(CO, A, B);
  specify
    specparam

      tplh$A$S  = 1.0,
      tphl$A$S  = 1.0,
      tplh$A$CO  = 1.0,
      tphl$A$CO  = 1.0,
      tplh$B$S  = 1.0,
      tphl$B$S  = 1.0,
      tplh$B$CO  = 1.0,
      tphl$B$CO  = 1.0;


     if (B == 1'b1)
	(A *> S) = (tplh$A$S,  tphl$A$S);
     if (B == 1'b0)
	(A *> S)  = (tplh$A$S,  tphl$A$S);
     if (A == 1'b1)
	(B *> S)  = (tplh$B$S,  tphl$B$S);
     if (A == 1'b0)
	(B *> S)  = (tplh$B$S,  tphl$B$S);
     (A *> CO) = (tplh$A$CO, tphl$A$CO);
     (B *> CO) = (tplh$B$CO, tphl$B$CO);

  endspecify
endmodule // ADDHX2MA10TR
`endcelldefine
//$Id: add.genpp,v 1.7 2006/06/01 15:56:41 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module ADDHX1P4MA10TR ( S, CO, A, B);
output S, CO;
input A, B;
  xor I0(S, A, B);
  and I1(CO, A, B);
  specify
    specparam

      tplh$A$S  = 1.0,
      tphl$A$S  = 1.0,
      tplh$A$CO  = 1.0,
      tphl$A$CO  = 1.0,
      tplh$B$S  = 1.0,
      tphl$B$S  = 1.0,
      tplh$B$CO  = 1.0,
      tphl$B$CO  = 1.0;


     if (B == 1'b1)
	(A *> S) = (tplh$A$S,  tphl$A$S);
     if (B == 1'b0)
	(A *> S)  = (tplh$A$S,  tphl$A$S);
     if (A == 1'b1)
	(B *> S)  = (tplh$B$S,  tphl$B$S);
     if (A == 1'b0)
	(B *> S)  = (tplh$B$S,  tphl$B$S);
     (A *> CO) = (tplh$A$CO, tphl$A$CO);
     (B *> CO) = (tplh$B$CO, tphl$B$CO);

  endspecify
endmodule // ADDHX1P4MA10TR
`endcelldefine
//$Id: add.genpp,v 1.7 2006/06/01 15:56:41 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module ADDHX1MA10TR ( S, CO, A, B);
output S, CO;
input A, B;
  xor I0(S, A, B);
  and I1(CO, A, B);
  specify
    specparam

      tplh$A$S  = 1.0,
      tphl$A$S  = 1.0,
      tplh$A$CO  = 1.0,
      tphl$A$CO  = 1.0,
      tplh$B$S  = 1.0,
      tphl$B$S  = 1.0,
      tplh$B$CO  = 1.0,
      tphl$B$CO  = 1.0;


     if (B == 1'b1)
	(A *> S) = (tplh$A$S,  tphl$A$S);
     if (B == 1'b0)
	(A *> S)  = (tplh$A$S,  tphl$A$S);
     if (A == 1'b1)
	(B *> S)  = (tplh$B$S,  tphl$B$S);
     if (A == 1'b0)
	(B *> S)  = (tplh$B$S,  tphl$B$S);
     (A *> CO) = (tplh$A$CO, tphl$A$CO);
     (B *> CO) = (tplh$B$CO, tphl$B$CO);

  endspecify
endmodule // ADDHX1MA10TR
`endcelldefine
//$Id: add.genpp,v 1.7 2006/06/01 15:56:41 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module ADDFX2MA10TR ( S, CO, A, B, CI);
output S, CO;
input A, B, CI;
  xor I0(S, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or  I4(CO, a_and_b, a_and_ci, b_and_ci);
  specify
    specparam

      tplh$A$S  = 1.0,
      tphl$A$S  = 1.0,
      tplh$A$CO  = 1.0,
      tphl$A$CO  = 1.0,
      tplh$B$S  = 1.0,
      tphl$B$S  = 1.0,
      tplh$B$CO  = 1.0,
      tphl$B$CO  = 1.0,
      tplh$CI$S  = 1.0,
      tphl$CI$S  = 1.0,
      tplh$CI$CO  = 1.0,
      tphl$CI$CO  = 1.0;


     if (B == 1'b0 && CI == 1'b0)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b1 && CI == 1'b1)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b0 && CI == 1'b1)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b1 && CI == 1'b0)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (A == 1'b0 && CI == 1'b0)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b1 && CI == 1'b1)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b0 && CI == 1'b1)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b1 && CI == 1'b0)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     
    if (B == 1'b1 && CI == 1'b0 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (B == 1'b0 && CI == 1'b1 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (A == 1'b1 && CI == 1'b0 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b0 && CI == 1'b1 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b1 && B == 1'b0 )
       (CI *> CO) = (tplh$CI$CO, tphl$CI$CO); 
    if (A == 1'b0 && B == 1'b1 )
       (CI *> CO) = (tplh$CI$CO, tphl$CI$CO); 
    if (A == 1'b0 && B == 1'b0 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S); 
    if (A == 1'b1 && B == 1'b1 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S); 
    if (A == 1'b0 && B == 1'b1 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S); 
    if (A == 1'b1 && B == 1'b0 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S);

  endspecify
endmodule // ADDFX2MA10TR
`endcelldefine
//$Id: add.genpp,v 1.7 2006/06/01 15:56:41 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module ADDFX1P4MA10TR ( S, CO, A, B, CI);
output S, CO;
input A, B, CI;
  xor I0(S, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or  I4(CO, a_and_b, a_and_ci, b_and_ci);
  specify
    specparam

      tplh$A$S  = 1.0,
      tphl$A$S  = 1.0,
      tplh$A$CO  = 1.0,
      tphl$A$CO  = 1.0,
      tplh$B$S  = 1.0,
      tphl$B$S  = 1.0,
      tplh$B$CO  = 1.0,
      tphl$B$CO  = 1.0,
      tplh$CI$S  = 1.0,
      tphl$CI$S  = 1.0,
      tplh$CI$CO  = 1.0,
      tphl$CI$CO  = 1.0;


     if (B == 1'b0 && CI == 1'b0)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b1 && CI == 1'b1)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b0 && CI == 1'b1)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b1 && CI == 1'b0)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (A == 1'b0 && CI == 1'b0)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b1 && CI == 1'b1)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b0 && CI == 1'b1)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b1 && CI == 1'b0)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     
    if (B == 1'b1 && CI == 1'b0 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (B == 1'b0 && CI == 1'b1 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (A == 1'b1 && CI == 1'b0 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b0 && CI == 1'b1 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b1 && B == 1'b0 )
       (CI *> CO) = (tplh$CI$CO, tphl$CI$CO); 
    if (A == 1'b0 && B == 1'b1 )
       (CI *> CO) = (tplh$CI$CO, tphl$CI$CO); 
    if (A == 1'b0 && B == 1'b0 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S); 
    if (A == 1'b1 && B == 1'b1 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S); 
    if (A == 1'b0 && B == 1'b1 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S); 
    if (A == 1'b1 && B == 1'b0 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S);

  endspecify
endmodule // ADDFX1P4MA10TR
`endcelldefine
//$Id: add.genpp,v 1.7 2006/06/01 15:56:41 kvaz Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module ADDFX1MA10TR ( S, CO, A, B, CI);
output S, CO;
input A, B, CI;
  xor I0(S, A, B, CI);
  and I1(a_and_b, A, B);
  and I2(a_and_ci, A, CI);
  and I3(b_and_ci, B, CI);
  or  I4(CO, a_and_b, a_and_ci, b_and_ci);
  specify
    specparam

      tplh$A$S  = 1.0,
      tphl$A$S  = 1.0,
      tplh$A$CO  = 1.0,
      tphl$A$CO  = 1.0,
      tplh$B$S  = 1.0,
      tphl$B$S  = 1.0,
      tplh$B$CO  = 1.0,
      tphl$B$CO  = 1.0,
      tplh$CI$S  = 1.0,
      tphl$CI$S  = 1.0,
      tplh$CI$CO  = 1.0,
      tphl$CI$CO  = 1.0;


     if (B == 1'b0 && CI == 1'b0)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b1 && CI == 1'b1)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b0 && CI == 1'b1)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (B == 1'b1 && CI == 1'b0)
	(A  *> S)  = (tplh$A$S,   tphl$A$S);
     if (A == 1'b0 && CI == 1'b0)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b1 && CI == 1'b1)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b0 && CI == 1'b1)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     if (A == 1'b1 && CI == 1'b0)
	(B  *> S)  = (tplh$B$S,   tphl$B$S);
     
    if (B == 1'b1 && CI == 1'b0 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (B == 1'b0 && CI == 1'b1 )
       (A *> CO) = (tplh$A$CO, tphl$A$CO); 
    if (A == 1'b1 && CI == 1'b0 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b0 && CI == 1'b1 )
       (B *> CO) = (tplh$B$CO, tphl$B$CO); 
    if (A == 1'b1 && B == 1'b0 )
       (CI *> CO) = (tplh$CI$CO, tphl$CI$CO); 
    if (A == 1'b0 && B == 1'b1 )
       (CI *> CO) = (tplh$CI$CO, tphl$CI$CO); 
    if (A == 1'b0 && B == 1'b0 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S); 
    if (A == 1'b1 && B == 1'b1 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S); 
    if (A == 1'b0 && B == 1'b1 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S); 
    if (A == 1'b1 && B == 1'b0 )
       (CI *> S) = (tplh$CI$S, tphl$CI$S);

  endspecify
endmodule // ADDFX1MA10TR
`endcelldefine
//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module A2SDFFQNX3MA10TR (QN, A, B, SI, SE, CK);
output QN;
input A, B, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  and     I0 (n2, A, B);
  udp_mux I2 (n1, n2, SI, SE);
  udp_dff I1 (n0, n1, clk, xRN, xSN, NOTIFIER);
  not     I3 (QN, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  and     I30 (SandRandSEbandB, B, SandRandSEb);
  and     I31 (SandRandSEbandA, A, SandRandSEb);
  specify
    specparam 
      tplh$CK$QN = 1.0,
      tphl$CK$QN = 1.0,
      tsetup$A$CK = 1.0,
      thold$A$CK = 0.5,
      tsetup$B$CK = 1.0,
      thold$B$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEbandB )
      (posedge CK *> (QN    -: A)) = (tplh$CK$QN,    tphl$CK$QN);
    if ( SandRandSEbandA )
      (posedge CK *> (QN    -: B)) = (tplh$CK$QN,    tphl$CK$QN);
    if ( SandRandSE )
      (posedge CK *> (QN    -: SI)) = (tplh$CK$QN,    tphl$CK$QN);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge A, tsetup$A$CK  ,thold$A$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge A, tsetup$A$CK  ,thold$A$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge B, tsetup$B$CK  ,thold$B$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge B, tsetup$B$CK  ,thold$B$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // A2SDFFQNX3MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module A2SDFFQNX2MA10TR (QN, A, B, SI, SE, CK);
output QN;
input A, B, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  and     I0 (n2, A, B);
  udp_mux I2 (n1, n2, SI, SE);
  udp_dff I1 (n0, n1, clk, xRN, xSN, NOTIFIER);
  not     I3 (QN, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  and     I30 (SandRandSEbandB, B, SandRandSEb);
  and     I31 (SandRandSEbandA, A, SandRandSEb);
  specify
    specparam 
      tplh$CK$QN = 1.0,
      tphl$CK$QN = 1.0,
      tsetup$A$CK = 1.0,
      thold$A$CK = 0.5,
      tsetup$B$CK = 1.0,
      thold$B$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEbandB )
      (posedge CK *> (QN    -: A)) = (tplh$CK$QN,    tphl$CK$QN);
    if ( SandRandSEbandA )
      (posedge CK *> (QN    -: B)) = (tplh$CK$QN,    tphl$CK$QN);
    if ( SandRandSE )
      (posedge CK *> (QN    -: SI)) = (tplh$CK$QN,    tphl$CK$QN);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge A, tsetup$A$CK  ,thold$A$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge A, tsetup$A$CK  ,thold$A$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge B, tsetup$B$CK  ,thold$B$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge B, tsetup$B$CK  ,thold$B$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // A2SDFFQNX2MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module A2SDFFQNX1MA10TR (QN, A, B, SI, SE, CK);
output QN;
input A, B, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  and     I0 (n2, A, B);
  udp_mux I2 (n1, n2, SI, SE);
  udp_dff I1 (n0, n1, clk, xRN, xSN, NOTIFIER);
  not     I3 (QN, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  and     I30 (SandRandSEbandB, B, SandRandSEb);
  and     I31 (SandRandSEbandA, A, SandRandSEb);
  specify
    specparam 
      tplh$CK$QN = 1.0,
      tphl$CK$QN = 1.0,
      tsetup$A$CK = 1.0,
      thold$A$CK = 0.5,
      tsetup$B$CK = 1.0,
      thold$B$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEbandB )
      (posedge CK *> (QN    -: A)) = (tplh$CK$QN,    tphl$CK$QN);
    if ( SandRandSEbandA )
      (posedge CK *> (QN    -: B)) = (tplh$CK$QN,    tphl$CK$QN);
    if ( SandRandSE )
      (posedge CK *> (QN    -: SI)) = (tplh$CK$QN,    tphl$CK$QN);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge A, tsetup$A$CK  ,thold$A$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge A, tsetup$A$CK  ,thold$A$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge B, tsetup$B$CK  ,thold$B$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge B, tsetup$B$CK  ,thold$B$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // A2SDFFQNX1MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module A2SDFFQNX0P5MA10TR (QN, A, B, SI, SE, CK);
output QN;
input A, B, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  and     I0 (n2, A, B);
  udp_mux I2 (n1, n2, SI, SE);
  udp_dff I1 (n0, n1, clk, xRN, xSN, NOTIFIER);
  not     I3 (QN, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  and     I30 (SandRandSEbandB, B, SandRandSEb);
  and     I31 (SandRandSEbandA, A, SandRandSEb);
  specify
    specparam 
      tplh$CK$QN = 1.0,
      tphl$CK$QN = 1.0,
      tsetup$A$CK = 1.0,
      thold$A$CK = 0.5,
      tsetup$B$CK = 1.0,
      thold$B$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEbandB )
      (posedge CK *> (QN    -: A)) = (tplh$CK$QN,    tphl$CK$QN);
    if ( SandRandSEbandA )
      (posedge CK *> (QN    -: B)) = (tplh$CK$QN,    tphl$CK$QN);
    if ( SandRandSE )
      (posedge CK *> (QN    -: SI)) = (tplh$CK$QN,    tphl$CK$QN);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge A, tsetup$A$CK  ,thold$A$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge A, tsetup$A$CK  ,thold$A$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge B, tsetup$B$CK  ,thold$B$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge B, tsetup$B$CK  ,thold$B$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // A2SDFFQNX0P5MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module A2SDFFQX4MA10TR (Q, A, B, SI, SE, CK);
output Q;
input A, B, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  and     I0 (n2, A, B);
  udp_mux I2 (n1, n2, SI, SE);
  udp_dff I1 (n0, n1, clk, xRN, xSN, NOTIFIER);
  buf     I3 (Q, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  and     I30 (SandRandSEbandB, B, SandRandSEb);
  and     I31 (SandRandSEbandA, A, SandRandSEb);
  specify
    specparam 
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$A$CK = 1.0,
      thold$A$CK = 0.5,
      tsetup$B$CK = 1.0,
      thold$B$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEbandB )
      (posedge CK *> (Q    +: A)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSEbandA )
      (posedge CK *> (Q    +: B)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge A, tsetup$A$CK  ,thold$A$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge A, tsetup$A$CK  ,thold$A$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge B, tsetup$B$CK  ,thold$B$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge B, tsetup$B$CK  ,thold$B$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // A2SDFFQX4MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module A2SDFFQX3MA10TR (Q, A, B, SI, SE, CK);
output Q;
input A, B, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  and     I0 (n2, A, B);
  udp_mux I2 (n1, n2, SI, SE);
  udp_dff I1 (n0, n1, clk, xRN, xSN, NOTIFIER);
  buf     I3 (Q, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  and     I30 (SandRandSEbandB, B, SandRandSEb);
  and     I31 (SandRandSEbandA, A, SandRandSEb);
  specify
    specparam 
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$A$CK = 1.0,
      thold$A$CK = 0.5,
      tsetup$B$CK = 1.0,
      thold$B$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEbandB )
      (posedge CK *> (Q    +: A)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSEbandA )
      (posedge CK *> (Q    +: B)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge A, tsetup$A$CK  ,thold$A$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge A, tsetup$A$CK  ,thold$A$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge B, tsetup$B$CK  ,thold$B$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge B, tsetup$B$CK  ,thold$B$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // A2SDFFQX3MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module A2SDFFQX2MA10TR (Q, A, B, SI, SE, CK);
output Q;
input A, B, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  and     I0 (n2, A, B);
  udp_mux I2 (n1, n2, SI, SE);
  udp_dff I1 (n0, n1, clk, xRN, xSN, NOTIFIER);
  buf     I3 (Q, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  and     I30 (SandRandSEbandB, B, SandRandSEb);
  and     I31 (SandRandSEbandA, A, SandRandSEb);
  specify
    specparam 
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$A$CK = 1.0,
      thold$A$CK = 0.5,
      tsetup$B$CK = 1.0,
      thold$B$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEbandB )
      (posedge CK *> (Q    +: A)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSEbandA )
      (posedge CK *> (Q    +: B)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge A, tsetup$A$CK  ,thold$A$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge A, tsetup$A$CK  ,thold$A$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge B, tsetup$B$CK  ,thold$B$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge B, tsetup$B$CK  ,thold$B$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // A2SDFFQX2MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module A2SDFFQX1MA10TR (Q, A, B, SI, SE, CK);
output Q;
input A, B, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  and     I0 (n2, A, B);
  udp_mux I2 (n1, n2, SI, SE);
  udp_dff I1 (n0, n1, clk, xRN, xSN, NOTIFIER);
  buf     I3 (Q, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  and     I30 (SandRandSEbandB, B, SandRandSEb);
  and     I31 (SandRandSEbandA, A, SandRandSEb);
  specify
    specparam 
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$A$CK = 1.0,
      thold$A$CK = 0.5,
      tsetup$B$CK = 1.0,
      thold$B$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEbandB )
      (posedge CK *> (Q    +: A)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSEbandA )
      (posedge CK *> (Q    +: B)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge A, tsetup$A$CK  ,thold$A$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge A, tsetup$A$CK  ,thold$A$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge B, tsetup$B$CK  ,thold$B$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge B, tsetup$B$CK  ,thold$B$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // A2SDFFQX1MA10TR
`endcelldefine
	

//$Id: sdff.genpp,v 1.18 2006/07/13 05:44:25 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module A2SDFFQX0P5MA10TR (Q, A, B, SI, SE, CK);
output Q;
input A, B, SI, SE, CK;
reg NOTIFIER;
supply1 xRN, xSN;
supply1 dRN, dSN;
  buf     IC (clk, CK);
  and     I0 (n2, A, B);
  udp_mux I2 (n1, n2, SI, SE);
  udp_dff I1 (n0, n1, clk, xRN, xSN, NOTIFIER);
  buf     I3 (Q, n0);
  and     I4 (SandR, xSN, xRN);
  and     I5 (SandRandSE, SandR, SE);
  not     I6 (SEb, SE);
  and     I7 (SandRandSEb, SandR, SEb);
  and     I30 (SandRandSEbandB, B, SandRandSEb);
  and     I31 (SandRandSEbandA, A, SandRandSEb);
  specify
    specparam 
      tplh$CK$Q = 1.0,
      tphl$CK$Q = 1.0,
      tsetup$A$CK = 1.0,
      thold$A$CK = 0.5,
      tsetup$B$CK = 1.0,
      thold$B$CK = 0.5,
      tsetup$SI$CK = 1.0,
      thold$SI$CK = 0.5,
      tsetup$SE$CK = 1.0,
      thold$SE$CK = 0.5,
      tminpwl$CK = 1.0,
      tminpwh$CK = 1.0,
      tperiod$CK = 1.0;
 // path delays
    if ( SandRandSEbandB )
      (posedge CK *> (Q    +: A)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSEbandA )
      (posedge CK *> (Q    +: B)) = (tplh$CK$Q,    tphl$CK$Q);
    if ( SandRandSE )
      (posedge CK *> (Q    +: SI)) = (tplh$CK$Q,    tphl$CK$Q);

// timing checks
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge A, tsetup$A$CK  ,thold$A$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge A, tsetup$A$CK  ,thold$A$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), posedge B, tsetup$B$CK  ,thold$B$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSEb == 1), negedge B, tsetup$B$CK  ,thold$B$CK  , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), posedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandRandSE == 1), negedge SI, tsetup$SI$CK, thold$SI$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), posedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $setuphold(posedge CK &&& (SandR == 1), negedge SE, tsetup$SE$CK, thold$SE$CK , NOTIFIER);
    $width(negedge CK &&& (SandR == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (SandR == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (SandR == 1), tperiod$CK, NOTIFIER);

endspecify
endmodule // A2SDFFQX0P5MA10TR
`endcelldefine
	

//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module A2DFFQNX3MA10TR (QN, A, B, CK);
output QN;
input  A, B, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  and     IA (n1, A, B);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  and     I30 (flagA, flag, B);
  and     I31 (flagB, flag, A);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$CK$QN	= 1.0,
    tphl$CK$QN	= 1.0,
    tsetup$A$CK	= 1.0,
    thold$A$CK	= 0.5,
    tsetup$B$CK	= 1.0,
    thold$B$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;

    if (flagA)
      (posedge CK *> (QN -: A)) = (tplh$CK$QN,   tphl$CK$QN);
    if (flagB)
      (posedge CK *> (QN -: B)) = (tplh$CK$QN,   tphl$CK$QN);
    $setuphold(posedge CK &&& (flag == 1), posedge A, tsetup$A$CK, thold$A$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge A, tsetup$A$CK, thold$A$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), posedge B, tsetup$B$CK, thold$B$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge B, tsetup$B$CK, thold$B$CK, NOTIFIER);
    $width(negedge CK &&& (flag  == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag  == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (flag  == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // A2DFFQNX3MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module A2DFFQNX2MA10TR (QN, A, B, CK);
output QN;
input  A, B, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  and     IA (n1, A, B);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  and     I30 (flagA, flag, B);
  and     I31 (flagB, flag, A);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$CK$QN	= 1.0,
    tphl$CK$QN	= 1.0,
    tsetup$A$CK	= 1.0,
    thold$A$CK	= 0.5,
    tsetup$B$CK	= 1.0,
    thold$B$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;

    if (flagA)
      (posedge CK *> (QN -: A)) = (tplh$CK$QN,   tphl$CK$QN);
    if (flagB)
      (posedge CK *> (QN -: B)) = (tplh$CK$QN,   tphl$CK$QN);
    $setuphold(posedge CK &&& (flag == 1), posedge A, tsetup$A$CK, thold$A$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge A, tsetup$A$CK, thold$A$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), posedge B, tsetup$B$CK, thold$B$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge B, tsetup$B$CK, thold$B$CK, NOTIFIER);
    $width(negedge CK &&& (flag  == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag  == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (flag  == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // A2DFFQNX2MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module A2DFFQNX1MA10TR (QN, A, B, CK);
output QN;
input  A, B, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  and     IA (n1, A, B);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  and     I30 (flagA, flag, B);
  and     I31 (flagB, flag, A);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$CK$QN	= 1.0,
    tphl$CK$QN	= 1.0,
    tsetup$A$CK	= 1.0,
    thold$A$CK	= 0.5,
    tsetup$B$CK	= 1.0,
    thold$B$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;

    if (flagA)
      (posedge CK *> (QN -: A)) = (tplh$CK$QN,   tphl$CK$QN);
    if (flagB)
      (posedge CK *> (QN -: B)) = (tplh$CK$QN,   tphl$CK$QN);
    $setuphold(posedge CK &&& (flag == 1), posedge A, tsetup$A$CK, thold$A$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge A, tsetup$A$CK, thold$A$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), posedge B, tsetup$B$CK, thold$B$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge B, tsetup$B$CK, thold$B$CK, NOTIFIER);
    $width(negedge CK &&& (flag  == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag  == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (flag  == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // A2DFFQNX1MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module A2DFFQNX0P5MA10TR (QN, A, B, CK);
output QN;
input  A, B, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  and     IA (n1, A, B);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  and     I30 (flagA, flag, B);
  and     I31 (flagB, flag, A);
  not     I2 (QN, n0);
  specify
    specparam
    tplh$CK$QN	= 1.0,
    tphl$CK$QN	= 1.0,
    tsetup$A$CK	= 1.0,
    thold$A$CK	= 0.5,
    tsetup$B$CK	= 1.0,
    thold$B$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;

    if (flagA)
      (posedge CK *> (QN -: A)) = (tplh$CK$QN,   tphl$CK$QN);
    if (flagB)
      (posedge CK *> (QN -: B)) = (tplh$CK$QN,   tphl$CK$QN);
    $setuphold(posedge CK &&& (flag == 1), posedge A, tsetup$A$CK, thold$A$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge A, tsetup$A$CK, thold$A$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), posedge B, tsetup$B$CK, thold$B$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge B, tsetup$B$CK, thold$B$CK, NOTIFIER);
    $width(negedge CK &&& (flag  == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag  == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (flag  == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // A2DFFQNX0P5MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module A2DFFQX4MA10TR (Q, A, B, CK);
output Q;
input  A, B, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  and     IA (n1, A, B);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  and     I30 (flagA, flag, B);
  and     I31 (flagB, flag, A);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$A$CK	= 1.0,
    thold$A$CK	= 0.5,
    tsetup$B$CK	= 1.0,
    thold$B$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;

    if (flagA)
      (posedge CK *> (Q +: A)) = (tplh$CK$Q,   tphl$CK$Q);
    if (flagB)
      (posedge CK *> (Q +: B)) = (tplh$CK$Q,   tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge A, tsetup$A$CK, thold$A$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge A, tsetup$A$CK, thold$A$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), posedge B, tsetup$B$CK, thold$B$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge B, tsetup$B$CK, thold$B$CK, NOTIFIER);
    $width(negedge CK &&& (flag  == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag  == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (flag  == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // A2DFFQX4MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module A2DFFQX3MA10TR (Q, A, B, CK);
output Q;
input  A, B, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  and     IA (n1, A, B);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  and     I30 (flagA, flag, B);
  and     I31 (flagB, flag, A);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$A$CK	= 1.0,
    thold$A$CK	= 0.5,
    tsetup$B$CK	= 1.0,
    thold$B$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;

    if (flagA)
      (posedge CK *> (Q +: A)) = (tplh$CK$Q,   tphl$CK$Q);
    if (flagB)
      (posedge CK *> (Q +: B)) = (tplh$CK$Q,   tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge A, tsetup$A$CK, thold$A$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge A, tsetup$A$CK, thold$A$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), posedge B, tsetup$B$CK, thold$B$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge B, tsetup$B$CK, thold$B$CK, NOTIFIER);
    $width(negedge CK &&& (flag  == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag  == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (flag  == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // A2DFFQX3MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module A2DFFQX2MA10TR (Q, A, B, CK);
output Q;
input  A, B, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  and     IA (n1, A, B);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  and     I30 (flagA, flag, B);
  and     I31 (flagB, flag, A);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$A$CK	= 1.0,
    thold$A$CK	= 0.5,
    tsetup$B$CK	= 1.0,
    thold$B$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;

    if (flagA)
      (posedge CK *> (Q +: A)) = (tplh$CK$Q,   tphl$CK$Q);
    if (flagB)
      (posedge CK *> (Q +: B)) = (tplh$CK$Q,   tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge A, tsetup$A$CK, thold$A$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge A, tsetup$A$CK, thold$A$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), posedge B, tsetup$B$CK, thold$B$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge B, tsetup$B$CK, thold$B$CK, NOTIFIER);
    $width(negedge CK &&& (flag  == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag  == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (flag  == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // A2DFFQX2MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module A2DFFQX1MA10TR (Q, A, B, CK);
output Q;
input  A, B, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  and     IA (n1, A, B);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  and     I30 (flagA, flag, B);
  and     I31 (flagB, flag, A);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$A$CK	= 1.0,
    thold$A$CK	= 0.5,
    tsetup$B$CK	= 1.0,
    thold$B$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;

    if (flagA)
      (posedge CK *> (Q +: A)) = (tplh$CK$Q,   tphl$CK$Q);
    if (flagB)
      (posedge CK *> (Q +: B)) = (tplh$CK$Q,   tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge A, tsetup$A$CK, thold$A$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge A, tsetup$A$CK, thold$A$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), posedge B, tsetup$B$CK, thold$B$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge B, tsetup$B$CK, thold$B$CK, NOTIFIER);
    $width(negedge CK &&& (flag  == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag  == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (flag  == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // A2DFFQX1MA10TR
`endcelldefine


//$Id: dff.genpp,v 1.15 2006/05/18 09:43:14 smd Exp $
//CONFIDENTIAL  AND  PROPRIETARY SOFTWARE OF ARM Physical IP, INC.
//
//Copyright (c) 1993-2006  ARM Physical IP, Inc.  All  Rights Reserved.
//
//Use of this Software is subject to the terms and conditions  of the
//applicable license agreement with ARM Physical IP, Inc.  In addition,
//this Software is protected by patents, copyright law and international
//treaties.
//
//The copyright notice(s) in this Software does not indicate actual or
//intended publication of this Software.
//

`timescale 1ns/1ps
`celldefine
module A2DFFQX0P5MA10TR (Q, A, B, CK);
output Q;
input  A, B, CK;
reg NOTIFIER;
supply1 xSN,xRN;
  buf     IC (clk, CK);
  and     IA (n1, A, B);
  udp_dff I0 (n0, n1, clk, xRN, xSN, NOTIFIER);
  and     I4 (flag, xRN, xSN);
  and     I30 (flagA, flag, B);
  and     I31 (flagB, flag, A);
  buf     I1 (Q, n0);
  specify
    specparam
    tplh$CK$Q	= 1.0,
    tphl$CK$Q	= 1.0,
    tsetup$A$CK	= 1.0,
    thold$A$CK	= 0.5,
    tsetup$B$CK	= 1.0,
    thold$B$CK	= 0.5,
    tminpwl$CK    = 1.0,
    tminpwh$CK    = 1.0,
    tperiod$CK    = 1.0;

    if (flagA)
      (posedge CK *> (Q +: A)) = (tplh$CK$Q,   tphl$CK$Q);
    if (flagB)
      (posedge CK *> (Q +: B)) = (tplh$CK$Q,   tphl$CK$Q);
    $setuphold(posedge CK &&& (flag == 1), posedge A, tsetup$A$CK, thold$A$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge A, tsetup$A$CK, thold$A$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), posedge B, tsetup$B$CK, thold$B$CK, NOTIFIER);
    $setuphold(posedge CK &&& (flag == 1), negedge B, tsetup$B$CK, thold$B$CK, NOTIFIER);
    $width(negedge CK &&& (flag  == 1), tminpwl$CK, 0, NOTIFIER);
    $width(posedge CK &&& (flag  == 1), tminpwh$CK, 0, NOTIFIER);
    $period(posedge CK &&& (flag  == 1), tperiod$CK, NOTIFIER);

   endspecify
endmodule // A2DFFQX0P5MA10TR
`endcelldefine



// This udp simulates the special latch behaviour of
// posticg cells.
primitive udp_plat (out, ena, ovrd, clock, NOTIFIER);
   output out;  
   input  ena, ovrd, clock, NOTIFIER;
   reg    out;

   table

// ovrd clock ena NOTIFIER : Qt : Qt+1
//
   1    ?    ?    ?   : ?  :  1  ;
   0    0    0    ?   : ?  :  0  ;
   0    0    1    ?   : ?  :  1  ;
   0    1    ?    ?   : ?  :  -  ;
   ?    1    *    ?   : ?  :  -  ; // no changes when in switches
   ?    ?    ?    *   : ?  :  x  ; // any notifier changed

   endtable
endprimitive // udp_plat


primitive udp_tlat (out, in, hold, clr_, set_, NOTIFIER);
   output out;  
   input  in, hold, clr_, set_, NOTIFIER;
   reg    out;

   table

// in  hold  clr_   set_  NOT  : Qt : Qt+1
//
   1  0   1   ?   ?   : ?  :  1  ; // 
   0  0   ?   1   ?   : ?  :  0  ; // 
   1  *   1   ?   ?   : 1  :  1  ; // reduce pessimism
   0  *   ?   1   ?   : 0  :  0  ; // reduce pessimism
   *  1   ?   ?   ?   : ?  :  -  ; // no changes when in switches
   ?  ?   ?   0   ?   : ?  :  1  ; // set output
   ?  1   1   *   ?   : 1  :  1  ; // cover all transistions on set_
   1  ?   1   *   ?   : 1  :  1  ; // cover all transistions on set_
   ?  ?   0   1   ?   : ?  :  0  ; // reset output
   ?  1   *   1   ?   : 0  :  0  ; // cover all transistions on clr_
   0  ?   *   1   ?   : 0  :  0  ; // cover all transistions on clr_
   ?  ?   ?   ?   *   : ?  :  x  ; // any notifier changed

   endtable
endprimitive // udp_tlat

// This primitive table models the behaviour of
// a wired AND-OR function. There are 2 inputs
// with two enables.
// in1a and in2a are pins of And 'a'
// in1b and in2b are pins of And 'b'
// out is an Or of And a and And b. 

primitive udp_wao (out, in1a, in1b, in2a, in2b);
   output out;
   input in1a, in1b, in2a, in2b;
  
   table

// in1a in1b in2a in2b: out
//
   1     1    1    ?  :  1;
   1     1    ?    1  :  1;
   0     0    1    ?  :  0;
   0     0    ?    1  :  0;
   1     ?    1    0  :  1;
   0     ?    1    0  :  0;
   ?     1    0    1  :  1;
   ?     0    0    1  :  0;

   endtable
endprimitive



primitive udp_sedff (out, in, clk, clr_, si, se, en, NOTIFIER);
   output out;  
   input  in, clk, clr_, si, se,  en, NOTIFIER;
   reg    out;

   table
   // in  clk  clr_  si  se  en  NOT : Qt : Qt+1
      ?    ?    ?     ?   ?   ?   *  : ?  :  x; // any notifier changed
      ?    ?    0     ?   ?   ?   ?  : ?  :  0;     
      ?    r    ?     0   1   ?   ?  : ?  :  0;     
      ?    r    1     1   1   ?   ?  : ?  :  1;
      ?    b    1     ?   *   ?   ?  : ?  :  -; // no changes when se switches
      ?    b    1     *   ?   ?   ?  : ?  :  -; // no changes when si switches
      *    b    1     ?   ?   ?   ?  : ?  :  -; // no changes when in switches
      *    ?    ?     ?   0   0   ?  : 0  :  0; // no changes when in switches
      ?    ?    ?     *   0   0   ?  : 0  :  0; // no changes when in switches
      ?    b    1     ?   ?   *   ?  : ?  :  -; // no changes when en switches
      ?    b    *     ?   ?   ?   ?  : 0  :  0; // no changes when en switches
      ?    ?    *     ?   0   0   ?  : 0  :  0; // no changes when en switches
      ?    b    ?     ?   ?   *   ?  : 0  :  0; // no changes when en switches
      ?    b    ?     ?   *   ?   ?  : 0  :  0; // no changes when en switches
      ?    b    ?     *   ?   ?   ?  : 0  :  0; // no changes when en switches
      *    b    ?     ?   ?   ?   ?  : 0  :  0; // no changes when en switches
      ?  (10)   ?     ?   ?   ?   ?  : ?  :  -;  // no changes on falling clk edge
      ?    *    1     1   1   ?   ?  : 1  :  1;
      ?    x    1     1   1   ?   ?  : 1  :  1;
      ?    *    1     1   ?   0   ?  : 1  :  1;
      ?    x    1     1   ?   0   ?  : 1  :  1;
      ?    *    ?     0   1   ?   ?  : 0  :  0;
      ?    x    ?     0   1   ?   ?  : 0  :  0;
      ?    *    ?     0   ?   0   ?  : 0  :  0;
      ?    x    ?     0   ?   0   ?  : 0  :  0;
      0    r    ?     0   ?   1   ?  : ?  :  0 ; 
      0    *    ?     0   ?   ?   ?  : 0  :  0 ; 
      0    x    ?     0   ?   ?   ?  : 0  :  0 ; 
      1    r    1     1   ?   1   ?  : ?  :  1 ; 
      1    *    1     1   ?   ?   ?  : 1  :  1 ; 
      1    x    1     1   ?   ?   ?  : 1  :  1 ; 
      ?  (x0)   ?     ?   ?   ?   ?  : ?  :  -;  // no changes on falling clk edge
      1    r    1     ?   0   1   ?  : ?  :  1;
      0    r    ?     ?   0   1   ?  : ?  :  0;
      ?    *    ?     ?   0   0   ?  : ?  :  -;
      ?    x    1     ?   0   0   ?  : ?  :  -;
      1    x    1     ?   0   ?   ?  : 1  :  1; // no changes when in switches
      0    x    ?     ?   0   ?   ?  : 0  :  0; // no changes when in switches
      1    x    ?     ?   0   0   ?  : 0  :  0; // no changes when in switches
      1    *    1     ?   0   ?   ?  : 1  :  1; // reduce pessimism
      0    *    ?     ?   0   ?   ?  : 0  :  0; // reduce pessimism

   endtable
endprimitive  /* udp_sedff */
   


primitive udp_mux (out, in, s_in, s_sel);
   output out;  
   input  in, s_in, s_sel;

   table

// in  s_in  s_sel :  out
//
   1  ?   0  :  1 ;
   0  ?   0  :  0 ;
   ?  1   1  :  1 ;
   ?  0   1  :  0 ;
   0  0   x  :  0 ;
   1  1   x  :  1 ;

   endtable
endprimitive // udp_mux


primitive udp_edff (out, in, clk, clr_, set_, en, NOTIFIER);
   output out;  
   input  in, clk, clr_, set_, en, NOTIFIER;
   reg    out;

   table

// in  clk  clr_   set_  en  NOT  : Qt : Qt+1
//
   0   r    ?      1     1   ?    : ?  :  0  ; // clock in 0
   1   r    1      ?     1   ?    : ?  :  1  ; // clock in 1
   ?   *    ?      ?     0   ?    : ?  :  -  ; // no changes, not enabled
   *   ?    ?      ?     0   ?    : ?  :  -  ; // no changes, not enabled
   1   *    1      ?     ?   ?    : 1  :  1  ; // reduce pessimism
   0   *    ?      1     ?   ?    : 0  :  0  ; // reduce pessimism
   ?   f    ?      ?     ?   ?    : ?  :  -  ; // no changes on negedge clk
   *   b    ?      ?     ?   ?    : ?  :  -  ; // no changes when in switches
   1   x    1      ?     ?   ?    : 1  :  1  ; // no changes when in switches
   0   x    ?      1     ?   ?    : 0  :  0  ; // no changes when in switches
   ?   b    ?      ?     *   ?    : ?  :  -  ; // no changes when en switches
   ?   x    1      1     0   ?    : ?  :  -  ; // no changes when en is disabled
   ?   ?    ?      0     ?   ?    : ?  :  1  ; // set output
   ?   b    1      *     ?   ?    : 1  :  1  ; // cover all transistions on set_
   ?   ?    1      *     0   ?    : 1  :  1  ; // cover all transistions on set_
   ?   ?    0      1     ?   ?    : ?  :  0  ; // reset output
   ?   b    *      1     ?   ?    : 0  :  0  ; // cover all transistions on clr_
   ?   ?    *      1     0   ?    : 0  :  0  ; // cover all transistions on clr_
   ?   ?    ?      ?     ?   *    : ?  :  x  ; // any notifier changed

   endtable
endprimitive // udp_edff


primitive udp_outrf (out, in, rwn, rw);
   output out;  
   input  in, rwn, rw;

   table

// in  rwn   rw   : out;
//	     	  
   0   0     ?    : 1  ; // 
   1   ?     1    : 1  ; // 
   ?   1     0    : 0  ; // 
   1   ?     0    : 0  ; // 
   0   1     ?    : 0  ; // 

   endtable
endprimitive // udp_outrf



primitive udp_dff (out, in, clk, clr_, set_, NOTIFIER);
   output out;  
   input  in, clk, clr_, set_, NOTIFIER;
   reg    out;

   table

// in  clk  clr_   set_  NOT  : Qt : Qt+1
//
   0  r   ?   1   ?   : ?  :  0  ; // clock in 0
   1  r   1   ?   ?   : ?  :  1  ; // clock in 1
   1  *   1   ?   ?   : 1  :  1  ; // reduce pessimism
   0  *   ?   1   ?   : 0  :  0  ; // reduce pessimism
   ?  f   ?   ?   ?   : ?  :  -  ; // no changes on negedge clk
   *  b   ?   ?   ?   : ?  :  -  ; // no changes when in switches
   ?  ?   ?   0   ?   : ?  :  1  ; // set output
   ?  b   1   *   ?   : 1  :  1  ; // cover all transistions on set_
   1  x   1   *   ?   : 1  :  1  ; // cover all transistions on set_
   ?  ?   0   1   ?   : ?  :  0  ; // reset output
   ?  b   *   1   ?   : 0  :  0  ; // cover all transistions on clr_
   0  x   *   1   ?   : 0  :  0  ; // cover all transistions on clr_
   ?  ?   ?   ?   *   : ?  :  x  ; // any notifier changed

   endtable
endprimitive // udp_dff


primitive udp_mux2 (out, in0, in1, sel);
   output out;  
   input  in0, in1, sel;

   table

// in0 in1  sel :  out
//
   1  ?   0  :  1 ;
   0  ?   0  :  0 ;
   ?  1   1  :  1 ;
   ?  0   1  :  0 ;
   0  0   x  :  0 ;
   1  1   x  :  1 ;

   endtable
endprimitive // udp_mux2


primitive udp_tlatrf (out, in, ww, wwn, NOTIFIER);
   output out;  
   input  in, ww, wwn, NOTIFIER;
   reg    out;

   table

// in  ww    wwn  NOT  : Qt : Qt+1
//	     
   1   ?     0    ?    : ?  :  1  ; // 
   1   1     ?    ?    : ?  :  1  ; // 
   0   ?     0    ?    : ?  :  0  ; // 
   0   1     ?    ?    : ?  :  0  ; // 
   1   *     ?    ?    : 1  :  1  ; // reduce pessimism
   1   ?     *    ?    : 1  :  1  ; // reduce pessimism
   0   *     ?    ?    : 0  :  0  ; // reduce pessimism
   0   ?     *    ?    : 0  :  0  ; // reduce pessimism
   *   0     1    ?    : ?  :  -  ; // no changes when in switches
   ?   ?     ?    *    : ?  :  x  ; // any notifier changed

   endtable
endprimitive // udp_tlatrf



primitive udp_mux4 (out, in0, in1, in2, in3, sel_0, sel_1);
   output out;  
   input  in0, in1, in2, in3, sel_0, sel_1;

   table

// in0 in1 in2 in3 sel_0 sel_1 :  out
//
   0  ?  ?  ?  0  0  :  0;
   1  ?  ?  ?  0  0  :  1;
   ?  0  ?  ?  1  0  :  0;
   ?  1  ?  ?  1  0  :  1;
   ?  ?  0  ?  0  1  :  0;
   ?  ?  1  ?  0  1  :  1;
   ?  ?  ?  0  1  1  :  0;
   ?  ?  ?  1  1  1  :  1;
   0  0  ?  ?  x  0  :  0;
   1  1  ?  ?  x  0  :  1;
   ?  ?  0  0  x  1  :  0;
   ?  ?  1  1  x  1  :  1;
   0  ?  0  ?  0  x  :  0;
   1  ?  1  ?  0  x  :  1;
   ?  0  ?  0  1  x  :  0;
   ?  1  ?  1  1  x  :  1;
   1  1  1  1  x  x  :  1;
   0  0  0  0  x  x  :  0;

   endtable
endprimitive // udp_mux4
